module top();
wire wire_clk;
wire [8:0] wire_image_header;
wire [8:0] wire_num_images;
wire [7:0] wire_pixel_data;
wire wire_pixel_valid;
wire wire_reset;
wire wire_start;
wire [8:0] wire_count_image;
wire wire_finish_reordering;
wire wire_hash_calc_done;
wire wire_image_buffer_valid;
wire [8:0] wire_last_image;
wire wire_new_reference_is_done;
wire [8:0] wire_temp_new_reference;
wire   net1000;
wire   net1001;


specify
    specparam CDS_LIBNAME  = "testLib";
    specparam CDS_CELLNAME = "top";
    specparam CDS_VIEWNAME = "schematic";
endspecify

top_syn I0(.clk(wire_clk)
,.image_header(wire_image_header[8:0])
,.num_images(wire_num_images[8:0])
,.pixel_data(wire_pixel_data[7:0])
,.pixel_valid(wire_pixel_valid)
,.reset(wire_reset)
,.start(wire_start)
,.count_image(wire_count_image[8:0])
,.finish_reordering(wire_finish_reordering)
,.hash_calc_done(wire_hash_calc_done)
,.image_buffer_valid(wire_image_buffer_valid)
,.last_image(wire_last_image[8:0])
,.new_reference_is_done(wire_new_reference_is_done)
,.temp_new_reference(wire_temp_new_reference[8:0])
);

pv0a PAD_G1 ( );
pv0c PAD_G3 (.VSSC(VSS));
pvda PAD_I1 ( );
pvdc PAD_I3 (.VDDC(VDD));

pc3d01 I5 ( .CIN(wire_clk), .PAD(net100));
pc3d01 I6 ( .CIN(wire_image_header[8]), .PAD(net101));
pc3d01 I7 ( .CIN(wire_image_header[7]), .PAD(net102));
pc3d01 I8 ( .CIN(wire_image_header[6]), .PAD(net103));
pc3d01 I9 ( .CIN(wire_image_header[5]), .PAD(net104));
pc3d01 I10 ( .CIN(wire_image_header[4]), .PAD(net105));
pc3d01 I11 ( .CIN(wire_image_header[3]), .PAD(net106));
pc3d01 I12 ( .CIN(wire_image_header[2]), .PAD(net107));
pc3d01 I13 ( .CIN(wire_image_header[1]), .PAD(net108));
pc3d01 I14 ( .CIN(wire_image_header[0]), .PAD(net109));
pc3d01 I15 ( .CIN(wire_num_images[8]), .PAD(net110));
pc3d01 I16 ( .CIN(wire_num_images[7]), .PAD(net111));
pc3d01 I17 ( .CIN(wire_num_images[6]), .PAD(net112));
pc3d01 I18 ( .CIN(wire_num_images[5]), .PAD(net113));
pc3d01 I19 ( .CIN(wire_num_images[4]), .PAD(net114));
pc3d01 I20 ( .CIN(wire_num_images[3]), .PAD(net115));
pc3d01 I21 ( .CIN(wire_num_images[2]), .PAD(net116));
pc3d01 I22 ( .CIN(wire_num_images[1]), .PAD(net117));
pc3d01 I23 ( .CIN(wire_num_images[0]), .PAD(net118));
pc3d01 I24 ( .CIN(wire_pixel_data[7]), .PAD(net119));
pc3d01 I25 ( .CIN(wire_pixel_data[6]), .PAD(net120));
pc3d01 I26 ( .CIN(wire_pixel_data[5]), .PAD(net121));
pc3d01 I27 ( .CIN(wire_pixel_data[4]), .PAD(net122));
pc3d01 I28 ( .CIN(wire_pixel_data[3]), .PAD(net123));
pc3d01 I29 ( .CIN(wire_pixel_data[2]), .PAD(net124));
pc3d01 I30 ( .CIN(wire_pixel_data[1]), .PAD(net125));
pc3d01 I31 ( .CIN(wire_pixel_data[0]), .PAD(net126));
pc3d01 I32 ( .CIN(wire_pixel_valid), .PAD(net127));
pc3d01 I33 ( .CIN(wire_reset), .PAD(net128));
pc3d01 I34 ( .CIN(wire_start), .PAD(net129));

pt3o01 I35 ( .PAD(net130), .I(wire_count_image[8]));
pt3o01 I36 ( .PAD(net131), .I(wire_count_image[7]));
pt3o01 I37 ( .PAD(net132), .I(wire_count_image[6]));
pt3o01 I38 ( .PAD(net133), .I(wire_count_image[5]));
pt3o01 I39 ( .PAD(net134), .I(wire_count_image[4]));
pt3o01 I40 ( .PAD(net135), .I(wire_count_image[3]));
pt3o01 I41 ( .PAD(net136), .I(wire_count_image[2]));
pt3o01 I42 ( .PAD(net137), .I(wire_count_image[1]));
pt3o01 I43 ( .PAD(net138), .I(wire_count_image[0]));
pt3o01 I44 ( .PAD(net139), .I(wire_finish_reordering));
pt3o01 I45 ( .PAD(net140), .I(wire_hash_calc_done));
pt3o01 I46 ( .PAD(net141), .I(wire_image_buffer_valid));
pt3o01 I47 ( .PAD(net142), .I(wire_last_image[8]));
pt3o01 I48 ( .PAD(net143), .I(wire_last_image[7]));
pt3o01 I49 ( .PAD(net144), .I(wire_last_image[6]));
pt3o01 I50 ( .PAD(net145), .I(wire_last_image[5]));
pt3o01 I51 ( .PAD(net146), .I(wire_last_image[4]));
pt3o01 I52 ( .PAD(net147), .I(wire_last_image[3]));
pt3o01 I53 ( .PAD(net148), .I(wire_last_image[2]));
pt3o01 I54 ( .PAD(net149), .I(wire_last_image[1]));
pt3o01 I55 ( .PAD(net150), .I(wire_last_image[0]));
pt3o01 I56 ( .PAD(net151), .I(wire_new_reference_is_done));
pt3o01 I57 ( .PAD(net152), .I(wire_temp_new_reference[8]));
pt3o01 I58 ( .PAD(net153), .I(wire_temp_new_reference[7]));
pt3o01 I59 ( .PAD(net154), .I(wire_temp_new_reference[6]));
pt3o01 I60 ( .PAD(net155), .I(wire_temp_new_reference[5]));
pt3o01 I61 ( .PAD(net156), .I(wire_temp_new_reference[4]));
pt3o01 I62 ( .PAD(net157), .I(wire_temp_new_reference[3]));
pt3o01 I63 ( .PAD(net158), .I(wire_temp_new_reference[2]));
pt3o01 I64 ( .PAD(net159), .I(wire_temp_new_reference[1]));
pt3o01 I65 ( .PAD(net160), .I(wire_temp_new_reference[0]));

pfrelr Pcornerlr();
pfrelr Pcornerll();
pfrelr Pcornerur();
pfrelr Pcornerul();

endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : U-2022.12
// Date      : Mon Feb 10 19:18:23 2025
/////////////////////////////////////////////////////////////


module image_buffer_DW01_inc_0_DW01_inc_5 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ah01d1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ah01d1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ah01d1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ah01d1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ah01d1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ah01d1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ah01d1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  inv0d0 U1 ( .I(A[0]), .ZN(SUM[0]) );
  xr02d1 U2 ( .A1(carry[8]), .A2(A[8]), .Z(SUM[8]) );
endmodule


module image_buffer ( clk, reset, pixel_data, pixel_valid, image_buffer_valid, 
        sum, buffer_I1, buffer_A1, buffer_WEB1 );
  input [7:0] pixel_data;
  output [15:0] sum;
  output [31:0] buffer_I1;
  output [11:0] buffer_A1;
  input clk, reset, pixel_valid;
  output image_buffer_valid, buffer_WEB1;
  wire   N13, N14, N15, N16, N17, N18, N19, N20, N21, N23, N24, N25, N26, N27,
         N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N51, N56, N57,
         N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N85, n10, n11, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90,
         N89, N88, N103, N102, N101, N100, \lte_52/A[5] , \lte_52/A[4] ,
         \add_38_aco/carry[15] , \add_38_aco/carry[14] ,
         \add_38_aco/carry[13] , \add_38_aco/carry[12] ,
         \add_38_aco/carry[11] , \add_38_aco/carry[10] , \add_38_aco/carry[9] ,
         \add_38_aco/carry[8] , \add_38_aco/carry[7] , \add_38_aco/carry[6] ,
         \add_38_aco/carry[5] , \add_38_aco/carry[4] , \add_38_aco/carry[3] ,
         \add_38_aco/carry[2] , \add_38_aco/carry[1] , n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62;
  wire   [8:0] pixel_index;
  assign buffer_WEB1 = 1'b0;
  assign buffer_I1[31] = 1'b0;
  assign buffer_I1[30] = 1'b0;
  assign buffer_I1[29] = 1'b0;
  assign buffer_I1[28] = 1'b0;
  assign buffer_I1[27] = 1'b0;
  assign buffer_I1[26] = 1'b0;
  assign buffer_I1[25] = 1'b0;
  assign buffer_I1[24] = 1'b0;
  assign buffer_I1[23] = 1'b0;
  assign buffer_I1[22] = 1'b0;
  assign buffer_I1[21] = 1'b0;
  assign buffer_I1[20] = 1'b0;
  assign buffer_I1[19] = 1'b0;
  assign buffer_I1[18] = 1'b0;
  assign buffer_I1[17] = 1'b0;
  assign buffer_I1[16] = 1'b0;
  assign buffer_I1[15] = 1'b0;
  assign buffer_I1[14] = 1'b0;
  assign buffer_I1[13] = 1'b0;
  assign buffer_I1[12] = 1'b0;
  assign buffer_I1[11] = 1'b0;
  assign buffer_I1[10] = 1'b0;
  assign buffer_I1[9] = 1'b0;
  assign buffer_I1[8] = 1'b0;

  dfcrn1 \pixel_index_reg[5]  ( .D(n39), .CP(clk), .CDN(n3), .QN(n11) );
  dfcrn1 \pixel_index_reg[4]  ( .D(n40), .CP(clk), .CDN(n3), .QN(n10) );
  lanhq1 \buffer_I1_reg[7]  ( .E(N51), .D(pixel_data[7]), .Q(buffer_I1[7]) );
  lanhq1 \buffer_I1_reg[6]  ( .E(N51), .D(pixel_data[6]), .Q(buffer_I1[6]) );
  lanhq1 \buffer_I1_reg[5]  ( .E(N51), .D(pixel_data[5]), .Q(buffer_I1[5]) );
  lanhq1 \buffer_I1_reg[4]  ( .E(N51), .D(pixel_data[4]), .Q(buffer_I1[4]) );
  lanhq1 \buffer_I1_reg[3]  ( .E(N51), .D(pixel_data[3]), .Q(buffer_I1[3]) );
  lanhq1 \buffer_I1_reg[2]  ( .E(N51), .D(pixel_data[2]), .Q(buffer_I1[2]) );
  lanhq1 \buffer_I1_reg[1]  ( .E(N51), .D(pixel_data[1]), .Q(buffer_I1[1]) );
  lanhq1 \buffer_I1_reg[0]  ( .E(N51), .D(pixel_data[0]), .Q(buffer_I1[0]) );
  lanhq1 \buffer_A1_reg[11]  ( .E(N51), .D(N74), .Q(buffer_A1[11]) );
  lanhq1 \buffer_A1_reg[10]  ( .E(N51), .D(N74), .Q(buffer_A1[10]) );
  lanhq1 \buffer_A1_reg[9]  ( .E(N51), .D(N74), .Q(buffer_A1[9]) );
  lanhq1 \buffer_A1_reg[8]  ( .E(N51), .D(N73), .Q(buffer_A1[8]) );
  lanhq1 \buffer_A1_reg[7]  ( .E(N51), .D(N72), .Q(buffer_A1[7]) );
  lanhq1 \buffer_A1_reg[6]  ( .E(N51), .D(N71), .Q(buffer_A1[6]) );
  lanhq1 \buffer_A1_reg[5]  ( .E(N51), .D(N70), .Q(buffer_A1[5]) );
  lanhq1 \buffer_A1_reg[4]  ( .E(N51), .D(N69), .Q(buffer_A1[4]) );
  lanhq1 \buffer_A1_reg[3]  ( .E(N51), .D(N68), .Q(buffer_A1[3]) );
  lanhq1 \buffer_A1_reg[2]  ( .E(N51), .D(N67), .Q(buffer_A1[2]) );
  lanhq1 \buffer_A1_reg[1]  ( .E(N51), .D(N66), .Q(buffer_A1[1]) );
  lanhq1 \buffer_A1_reg[0]  ( .E(N51), .D(N65), .Q(buffer_A1[0]) );
  image_buffer_DW01_inc_0_DW01_inc_5 add_33 ( .A({pixel_index[8:6], 
        \lte_52/A[5] , \lte_52/A[4] , pixel_index[3:0]}), .SUM({N21, N20, N19, 
        N18, N17, N16, N15, N14, N13}) );
  ad01d0 \add_38_aco/U1_1  ( .A(N89), .B(pixel_data[1]), .CI(
        \add_38_aco/carry[1] ), .CO(\add_38_aco/carry[2] ), .S(N24) );
  ad01d0 \add_38_aco/U1_2  ( .A(N90), .B(pixel_data[2]), .CI(
        \add_38_aco/carry[2] ), .CO(\add_38_aco/carry[3] ), .S(N25) );
  ad01d0 \add_38_aco/U1_3  ( .A(N91), .B(pixel_data[3]), .CI(
        \add_38_aco/carry[3] ), .CO(\add_38_aco/carry[4] ), .S(N26) );
  ad01d0 \add_38_aco/U1_4  ( .A(N92), .B(pixel_data[4]), .CI(
        \add_38_aco/carry[4] ), .CO(\add_38_aco/carry[5] ), .S(N27) );
  ad01d0 \add_38_aco/U1_5  ( .A(N93), .B(pixel_data[5]), .CI(
        \add_38_aco/carry[5] ), .CO(\add_38_aco/carry[6] ), .S(N28) );
  ad01d0 \add_38_aco/U1_6  ( .A(N94), .B(pixel_data[6]), .CI(
        \add_38_aco/carry[6] ), .CO(\add_38_aco/carry[7] ), .S(N29) );
  ad01d0 \add_38_aco/U1_7  ( .A(N95), .B(pixel_data[7]), .CI(
        \add_38_aco/carry[7] ), .CO(\add_38_aco/carry[8] ), .S(N30) );
  dfcrq1 image_buffer_valid_reg ( .D(n20), .CP(clk), .CDN(n3), .Q(
        image_buffer_valid) );
  dfcrq1 \sum_reg[15]  ( .D(n35), .CP(clk), .CDN(n1), .Q(sum[15]) );
  dfcrq1 \sum_reg[14]  ( .D(n34), .CP(clk), .CDN(n1), .Q(sum[14]) );
  dfcrq1 \sum_reg[13]  ( .D(n33), .CP(clk), .CDN(n2), .Q(sum[13]) );
  dfcrq1 \sum_reg[12]  ( .D(n32), .CP(clk), .CDN(n2), .Q(sum[12]) );
  dfcrq1 \sum_reg[11]  ( .D(n31), .CP(clk), .CDN(n2), .Q(sum[11]) );
  dfcrq1 \sum_reg[10]  ( .D(n30), .CP(clk), .CDN(n2), .Q(sum[10]) );
  dfcrq1 \sum_reg[9]  ( .D(n29), .CP(clk), .CDN(n2), .Q(sum[9]) );
  dfcrq1 \sum_reg[8]  ( .D(n28), .CP(clk), .CDN(n2), .Q(sum[8]) );
  dfcrq1 \sum_reg[7]  ( .D(n27), .CP(clk), .CDN(n2), .Q(sum[7]) );
  dfcrq1 \sum_reg[6]  ( .D(n26), .CP(clk), .CDN(n2), .Q(sum[6]) );
  dfcrq1 \sum_reg[5]  ( .D(n25), .CP(clk), .CDN(n2), .Q(sum[5]) );
  dfcrq1 \sum_reg[4]  ( .D(n24), .CP(clk), .CDN(n2), .Q(sum[4]) );
  dfcrq1 \sum_reg[3]  ( .D(n23), .CP(clk), .CDN(n3), .Q(sum[3]) );
  dfcrq1 \sum_reg[2]  ( .D(n22), .CP(clk), .CDN(n3), .Q(sum[2]) );
  dfcrq1 \sum_reg[1]  ( .D(n21), .CP(clk), .CDN(n3), .Q(sum[1]) );
  dfcrq1 \sum_reg[0]  ( .D(n36), .CP(clk), .CDN(n1), .Q(sum[0]) );
  dfcrq1 \pixel_index_reg[2]  ( .D(n42), .CP(clk), .CDN(n1), .Q(pixel_index[2]) );
  dfcrq1 \pixel_index_reg[7]  ( .D(n37), .CP(clk), .CDN(n1), .Q(pixel_index[7]) );
  dfcrq1 \pixel_index_reg[8]  ( .D(n44), .CP(clk), .CDN(n1), .Q(pixel_index[8]) );
  dfcrq1 \pixel_index_reg[6]  ( .D(n38), .CP(clk), .CDN(n1), .Q(pixel_index[6]) );
  dfcrq1 \pixel_index_reg[3]  ( .D(n41), .CP(clk), .CDN(n1), .Q(pixel_index[3]) );
  dfcrq1 \pixel_index_reg[0]  ( .D(n45), .CP(clk), .CDN(n1), .Q(pixel_index[0]) );
  dfcrq1 \pixel_index_reg[1]  ( .D(n43), .CP(clk), .CDN(n1), .Q(pixel_index[1]) );
  oan211d2 U6 ( .C1(n59), .C2(n60), .B(n19), .A(image_buffer_valid), .ZN(N51)
         );
  buffd1 U7 ( .I(N85), .Z(n4) );
  buffd1 U8 ( .I(N85), .Z(n6) );
  buffd1 U9 ( .I(N85), .Z(n5) );
  inv0d1 U31 ( .I(n19), .ZN(n54) );
  inv0d0 U32 ( .I(n14), .ZN(n16) );
  buffd1 U33 ( .I(n62), .Z(n2) );
  buffd1 U34 ( .I(n62), .Z(n1) );
  buffd1 U35 ( .I(n62), .Z(n3) );
  nd02d1 U36 ( .A1(pixel_valid), .A2(n46), .ZN(n19) );
  inv0d0 U37 ( .I(n15), .ZN(N63) );
  xr02d1 U38 ( .A1(\add_38_aco/carry[15] ), .A2(N103), .Z(N38) );
  an02d0 U39 ( .A1(N102), .A2(\add_38_aco/carry[14] ), .Z(
        \add_38_aco/carry[15] ) );
  xr02d1 U40 ( .A1(\add_38_aco/carry[14] ), .A2(N102), .Z(N37) );
  an02d0 U41 ( .A1(N101), .A2(\add_38_aco/carry[13] ), .Z(
        \add_38_aco/carry[14] ) );
  xr02d1 U42 ( .A1(\add_38_aco/carry[13] ), .A2(N101), .Z(N36) );
  an02d0 U43 ( .A1(N100), .A2(\add_38_aco/carry[12] ), .Z(
        \add_38_aco/carry[13] ) );
  xr02d1 U44 ( .A1(\add_38_aco/carry[12] ), .A2(N100), .Z(N35) );
  an02d0 U45 ( .A1(N99), .A2(\add_38_aco/carry[11] ), .Z(
        \add_38_aco/carry[12] ) );
  xr02d1 U46 ( .A1(\add_38_aco/carry[11] ), .A2(N99), .Z(N34) );
  an02d0 U47 ( .A1(N98), .A2(\add_38_aco/carry[10] ), .Z(
        \add_38_aco/carry[11] ) );
  xr02d1 U48 ( .A1(\add_38_aco/carry[10] ), .A2(N98), .Z(N33) );
  an02d0 U49 ( .A1(N97), .A2(\add_38_aco/carry[9] ), .Z(\add_38_aco/carry[10] ) );
  xr02d1 U50 ( .A1(\add_38_aco/carry[9] ), .A2(N97), .Z(N32) );
  an02d0 U51 ( .A1(N96), .A2(\add_38_aco/carry[8] ), .Z(\add_38_aco/carry[9] )
         );
  xr02d1 U52 ( .A1(\add_38_aco/carry[8] ), .A2(N96), .Z(N31) );
  an02d0 U53 ( .A1(N88), .A2(pixel_data[0]), .Z(\add_38_aco/carry[1] ) );
  xr02d1 U54 ( .A1(pixel_data[0]), .A2(N88), .Z(N23) );
  an02d0 U55 ( .A1(sum[0]), .A2(n4), .Z(N88) );
  an02d0 U56 ( .A1(sum[10]), .A2(n6), .Z(N98) );
  an02d0 U57 ( .A1(sum[11]), .A2(n6), .Z(N99) );
  an02d0 U58 ( .A1(sum[12]), .A2(n6), .Z(N100) );
  an02d0 U59 ( .A1(sum[13]), .A2(n6), .Z(N101) );
  an02d0 U60 ( .A1(sum[14]), .A2(n6), .Z(N102) );
  an02d0 U61 ( .A1(sum[15]), .A2(n5), .Z(N103) );
  an02d0 U62 ( .A1(sum[1]), .A2(n6), .Z(N89) );
  an02d0 U63 ( .A1(sum[2]), .A2(n6), .Z(N90) );
  an02d0 U64 ( .A1(sum[3]), .A2(n5), .Z(N91) );
  an02d0 U65 ( .A1(sum[4]), .A2(n5), .Z(N92) );
  an02d0 U66 ( .A1(sum[5]), .A2(n5), .Z(N93) );
  an02d0 U67 ( .A1(sum[6]), .A2(n5), .Z(N94) );
  an02d0 U68 ( .A1(sum[7]), .A2(n5), .Z(N95) );
  an02d0 U69 ( .A1(sum[8]), .A2(n5), .Z(N96) );
  an02d0 U70 ( .A1(n6), .A2(sum[9]), .Z(N97) );
  nd12d0 U71 ( .A1(pixel_index[1]), .A2(n17), .ZN(n7) );
  oaim21d1 U72 ( .B1(pixel_index[0]), .B2(pixel_index[1]), .A(n7), .ZN(N56) );
  or02d0 U73 ( .A1(n7), .A2(pixel_index[2]), .Z(n8) );
  oaim21d1 U74 ( .B1(n7), .B2(pixel_index[2]), .A(n8), .ZN(N57) );
  or02d0 U75 ( .A1(n8), .A2(pixel_index[3]), .Z(n9) );
  oaim21d1 U76 ( .B1(n8), .B2(pixel_index[3]), .A(n9), .ZN(N58) );
  or02d0 U77 ( .A1(n9), .A2(\lte_52/A[4] ), .Z(n12) );
  oaim21d1 U78 ( .B1(n9), .B2(\lte_52/A[4] ), .A(n12), .ZN(N59) );
  or02d0 U79 ( .A1(n12), .A2(\lte_52/A[5] ), .Z(n13) );
  oaim21d1 U80 ( .B1(n12), .B2(\lte_52/A[5] ), .A(n13), .ZN(N60) );
  nr02d0 U81 ( .A1(n13), .A2(pixel_index[6]), .ZN(n14) );
  oaim21d1 U82 ( .B1(n13), .B2(pixel_index[6]), .A(n16), .ZN(N61) );
  xr02d1 U83 ( .A1(pixel_index[7]), .A2(n14), .Z(N62) );
  nr03d0 U84 ( .A1(pixel_index[7]), .A2(pixel_index[8]), .A3(n16), .ZN(N64) );
  oan211d1 U85 ( .C1(n16), .C2(pixel_index[7]), .B(pixel_index[8]), .A(N64), 
        .ZN(n15) );
  inv0d0 U86 ( .I(reset), .ZN(n62) );
  oai22d1 U87 ( .A1(pixel_valid), .A2(n17), .B1(n18), .B2(n19), .ZN(n45) );
  inv0d0 U88 ( .I(N13), .ZN(n18) );
  oai22d1 U89 ( .A1(pixel_valid), .A2(n46), .B1(n47), .B2(n19), .ZN(n44) );
  inv0d0 U90 ( .I(N21), .ZN(n47) );
  oai22d1 U91 ( .A1(pixel_valid), .A2(n48), .B1(n49), .B2(n19), .ZN(n43) );
  inv0d0 U92 ( .I(N14), .ZN(n49) );
  inv0d0 U93 ( .I(pixel_index[1]), .ZN(n48) );
  oai22d1 U94 ( .A1(pixel_valid), .A2(n50), .B1(n51), .B2(n19), .ZN(n42) );
  inv0d0 U95 ( .I(N15), .ZN(n51) );
  oai22d1 U96 ( .A1(pixel_valid), .A2(n52), .B1(n53), .B2(n19), .ZN(n41) );
  inv0d0 U97 ( .I(N16), .ZN(n53) );
  oaim22d1 U98 ( .A1(pixel_valid), .A2(n10), .B1(N17), .B2(n54), .ZN(n40) );
  oaim22d1 U99 ( .A1(pixel_valid), .A2(n11), .B1(N18), .B2(n54), .ZN(n39) );
  oaim22d1 U100 ( .A1(pixel_valid), .A2(n55), .B1(N19), .B2(n54), .ZN(n38) );
  oaim22d1 U101 ( .A1(pixel_valid), .A2(n56), .B1(N20), .B2(n54), .ZN(n37) );
  mx02d1 U102 ( .I0(N23), .I1(sum[0]), .S(n19), .Z(n36) );
  mx02d1 U103 ( .I0(N38), .I1(sum[15]), .S(n19), .Z(n35) );
  mx02d1 U104 ( .I0(N37), .I1(sum[14]), .S(n19), .Z(n34) );
  mx02d1 U105 ( .I0(sum[13]), .I1(N36), .S(n54), .Z(n33) );
  mx02d1 U106 ( .I0(sum[12]), .I1(N35), .S(n54), .Z(n32) );
  mx02d1 U107 ( .I0(sum[11]), .I1(N34), .S(n54), .Z(n31) );
  mx02d1 U108 ( .I0(sum[10]), .I1(N33), .S(n54), .Z(n30) );
  mx02d1 U109 ( .I0(sum[9]), .I1(N32), .S(n54), .Z(n29) );
  mx02d1 U110 ( .I0(sum[8]), .I1(N31), .S(n54), .Z(n28) );
  mx02d1 U111 ( .I0(sum[7]), .I1(N30), .S(n54), .Z(n27) );
  mx02d1 U112 ( .I0(sum[6]), .I1(N29), .S(n54), .Z(n26) );
  mx02d1 U113 ( .I0(sum[5]), .I1(N28), .S(n54), .Z(n25) );
  mx02d1 U114 ( .I0(sum[4]), .I1(N27), .S(n54), .Z(n24) );
  mx02d1 U115 ( .I0(sum[3]), .I1(N26), .S(n54), .Z(n23) );
  mx02d1 U116 ( .I0(sum[2]), .I1(N25), .S(n54), .Z(n22) );
  mx02d1 U117 ( .I0(sum[1]), .I1(N24), .S(n54), .Z(n21) );
  mx02d1 U118 ( .I0(image_buffer_valid), .I1(pixel_index[8]), .S(pixel_valid), 
        .Z(n20) );
  an02d0 U119 ( .A1(N64), .A2(n5), .Z(N74) );
  an02d0 U120 ( .A1(N63), .A2(n4), .Z(N73) );
  an02d0 U121 ( .A1(N62), .A2(n4), .Z(N72) );
  an02d0 U122 ( .A1(N61), .A2(n4), .Z(N71) );
  an02d0 U123 ( .A1(N60), .A2(n4), .Z(N70) );
  an02d0 U124 ( .A1(N59), .A2(n4), .Z(N69) );
  an02d0 U125 ( .A1(N58), .A2(n4), .Z(N68) );
  an02d0 U126 ( .A1(N57), .A2(n4), .Z(N67) );
  an02d0 U127 ( .A1(N56), .A2(n4), .Z(N66) );
  an02d0 U128 ( .A1(n17), .A2(n5), .Z(N65) );
  nd04d0 U129 ( .A1(n50), .A2(n52), .A3(n57), .A4(n58), .ZN(N85) );
  nr04d0 U130 ( .A1(pixel_index[1]), .A2(pixel_index[0]), .A3(\lte_52/A[5] ), 
        .A4(\lte_52/A[4] ), .ZN(n58) );
  inv0d0 U131 ( .I(n10), .ZN(\lte_52/A[4] ) );
  inv0d0 U132 ( .I(n11), .ZN(\lte_52/A[5] ) );
  nr03d0 U133 ( .A1(pixel_index[6]), .A2(pixel_index[8]), .A3(pixel_index[7]), 
        .ZN(n57) );
  inv0d0 U134 ( .I(pixel_index[2]), .ZN(n50) );
  inv0d0 U135 ( .I(pixel_index[8]), .ZN(n46) );
  nd04d0 U136 ( .A1(pixel_valid), .A2(n10), .A3(n11), .A4(n17), .ZN(n60) );
  inv0d0 U137 ( .I(pixel_index[0]), .ZN(n17) );
  nd04d0 U138 ( .A1(n55), .A2(n56), .A3(n52), .A4(n61), .ZN(n59) );
  nr02d0 U139 ( .A1(pixel_index[2]), .A2(pixel_index[1]), .ZN(n61) );
  inv0d0 U140 ( .I(pixel_index[3]), .ZN(n52) );
  inv0d0 U141 ( .I(pixel_index[7]), .ZN(n56) );
  inv0d0 U142 ( .I(pixel_index[6]), .ZN(n55) );
endmodule


module hash_calc_DW01_inc_1_DW01_inc_4 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ah01d1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ah01d1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ah01d1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ah01d1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ah01d1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ah01d1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ah01d1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  inv0d0 U1 ( .I(A[0]), .ZN(SUM[0]) );
  xr02d1 U2 ( .A1(carry[8]), .A2(A[8]), .Z(SUM[8]) );
endmodule


module hash_calc ( clk, reset, image_header, hash_start, sum, hash_calc_done, 
        hash_O2, hash_I1, hash_A1, hash_A2, hash_WEB1, hash_WEB2 );
  input [8:0] image_header;
  input [15:0] sum;
  input [31:0] hash_O2;
  output [31:0] hash_I1;
  output [11:0] hash_A1;
  output [11:0] hash_A2;
  input clk, reset, hash_start;
  output hash_calc_done, hash_WEB1, hash_WEB2;
  wire   bit_value, N149, N150, N151, N152, N153, N154, N155, N156, N157, N159,
         N160, N161, N162, N217, N218, N219, N220, N221, N222, N223, N224,
         N225, N226, N227, N228, N241, N242, N243, N244, N245, N246, N247,
         N248, N249, N250, N251, N252, N253, N254, N255, N256, N257, N258,
         N259, N260, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, n36, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         N203, N202, N201, N200, N199, N198, N197, N196, N195, N194, N193,
         N192, \add_49/carry[4] , \add_49/carry[3] , \add_49/carry[2] ,
         \add_0_root_add_0_root_sub_75/carry[11] ,
         \add_0_root_add_0_root_sub_75/carry[10] ,
         \add_0_root_add_0_root_sub_75/carry[9] ,
         \add_0_root_add_0_root_sub_75/carry[8] ,
         \add_0_root_add_0_root_sub_75/carry[7] ,
         \add_0_root_add_0_root_sub_75/carry[6] ,
         \add_0_root_add_0_root_sub_75/carry[5] ,
         \add_0_root_add_0_root_sub_75/carry[4] ,
         \add_0_root_add_0_root_sub_75/carry[3] ,
         \add_0_root_add_0_root_sub_75/carry[2] ,
         \add_1_root_add_0_root_sub_75/carry[11] ,
         \add_1_root_add_0_root_sub_75/carry[10] ,
         \add_1_root_add_0_root_sub_75/carry[9] ,
         \add_1_root_add_0_root_sub_75/carry[8] ,
         \add_1_root_add_0_root_sub_75/carry[7] ,
         \add_1_root_add_0_root_sub_75/carry[6] ,
         \add_1_root_add_0_root_sub_75/carry[5] ,
         \add_1_root_add_0_root_sub_75/carry[4] ,
         \add_1_root_add_0_root_sub_75/A[3] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n37, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231;
  assign hash_WEB1 = 1'b0;
  assign hash_A2[9] = 1'b0;
  assign hash_A2[10] = 1'b0;
  assign hash_A2[11] = 1'b0;
  assign hash_WEB2 = 1'b1;

  dfcrn1 \hash_index_reg[3]  ( .D(n186), .CP(clk), .CDN(n12), .QN(n36) );
  labhb1 \hash_A1_reg[11]  ( .E(n17), .D(N227), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[11]) );
  labhb1 \hash_A1_reg[10]  ( .E(n17), .D(N226), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[10]) );
  labhb1 \hash_A1_reg[9]  ( .E(n17), .D(N225), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[9]) );
  labhb1 \hash_A1_reg[8]  ( .E(n17), .D(N224), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[8]) );
  labhb1 \hash_A1_reg[7]  ( .E(n16), .D(N223), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[7]) );
  labhb1 \hash_A1_reg[6]  ( .E(n16), .D(N222), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[6]) );
  labhb1 \hash_A1_reg[5]  ( .E(n16), .D(N221), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[5]) );
  labhb1 \hash_A1_reg[4]  ( .E(n16), .D(N220), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[4]) );
  labhb1 \hash_A1_reg[3]  ( .E(n15), .D(N219), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[3]) );
  labhb1 \hash_A1_reg[2]  ( .E(n15), .D(N218), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[2]) );
  labhb1 \hash_A1_reg[1]  ( .E(n15), .D(N217), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[1]) );
  labhb1 \hash_A1_reg[0]  ( .E(n15), .D(n228), .CDN(1'b1), .SDN(n149), .Q(
        hash_A1[0]) );
  lanhq1 bit_value_reg ( .E(N273), .D(N274), .Q(bit_value) );
  dfcrn1 \bits_reg[31]  ( .D(n154), .CP(clk), .CDN(n12), .QN(n38) );
  lanhq1 \hash_I1_reg[31]  ( .E(n19), .D(N272), .Q(hash_I1[31]) );
  dfcrn1 \bits_reg[30]  ( .D(n155), .CP(clk), .CDN(n12), .QN(n39) );
  lanhq1 \hash_I1_reg[30]  ( .E(n19), .D(N271), .Q(hash_I1[30]) );
  dfcrn1 \bits_reg[29]  ( .D(n156), .CP(clk), .CDN(n12), .QN(n40) );
  lanhq1 \hash_I1_reg[29]  ( .E(n19), .D(N270), .Q(hash_I1[29]) );
  dfcrn1 \bits_reg[28]  ( .D(n157), .CP(clk), .CDN(n12), .QN(n41) );
  lanhq1 \hash_I1_reg[28]  ( .E(n19), .D(N269), .Q(hash_I1[28]) );
  dfcrn1 \bits_reg[27]  ( .D(n158), .CP(clk), .CDN(n12), .QN(n42) );
  lanhq1 \hash_I1_reg[27]  ( .E(n19), .D(N268), .Q(hash_I1[27]) );
  dfcrn1 \bits_reg[26]  ( .D(n159), .CP(clk), .CDN(n11), .QN(n43) );
  lanhq1 \hash_I1_reg[26]  ( .E(n19), .D(N267), .Q(hash_I1[26]) );
  dfcrn1 \bits_reg[25]  ( .D(n160), .CP(clk), .CDN(n11), .QN(n44) );
  lanhq1 \hash_I1_reg[25]  ( .E(n19), .D(N266), .Q(hash_I1[25]) );
  dfcrn1 \bits_reg[24]  ( .D(n161), .CP(clk), .CDN(n11), .QN(n45) );
  lanhq1 \hash_I1_reg[24]  ( .E(n19), .D(N265), .Q(hash_I1[24]) );
  dfcrn1 \bits_reg[23]  ( .D(n162), .CP(clk), .CDN(n11), .QN(n46) );
  lanhq1 \hash_I1_reg[23]  ( .E(n19), .D(N264), .Q(hash_I1[23]) );
  dfcrn1 \bits_reg[22]  ( .D(n163), .CP(clk), .CDN(n11), .QN(n47) );
  lanhq1 \hash_I1_reg[22]  ( .E(n20), .D(N263), .Q(hash_I1[22]) );
  dfcrn1 \bits_reg[21]  ( .D(n164), .CP(clk), .CDN(n11), .QN(n48) );
  lanhq1 \hash_I1_reg[21]  ( .E(n20), .D(N262), .Q(hash_I1[21]) );
  dfcrn1 \bits_reg[20]  ( .D(n165), .CP(clk), .CDN(n11), .QN(n49) );
  lanhq1 \hash_I1_reg[20]  ( .E(n20), .D(N261), .Q(hash_I1[20]) );
  dfcrn1 \bits_reg[19]  ( .D(n166), .CP(clk), .CDN(n11), .QN(n50) );
  lanhq1 \hash_I1_reg[19]  ( .E(n20), .D(N260), .Q(hash_I1[19]) );
  dfcrn1 \bits_reg[18]  ( .D(n167), .CP(clk), .CDN(n11), .QN(n51) );
  lanhq1 \hash_I1_reg[18]  ( .E(n20), .D(N259), .Q(hash_I1[18]) );
  dfcrn1 \bits_reg[17]  ( .D(n168), .CP(clk), .CDN(n11), .QN(n52) );
  lanhq1 \hash_I1_reg[17]  ( .E(n20), .D(N258), .Q(hash_I1[17]) );
  dfcrn1 \bits_reg[16]  ( .D(n169), .CP(clk), .CDN(n10), .QN(n53) );
  lanhq1 \hash_I1_reg[16]  ( .E(n20), .D(N257), .Q(hash_I1[16]) );
  dfcrn1 \bits_reg[15]  ( .D(n170), .CP(clk), .CDN(n10), .QN(n54) );
  lanhq1 \hash_I1_reg[15]  ( .E(n20), .D(N256), .Q(hash_I1[15]) );
  dfcrn1 \bits_reg[14]  ( .D(n171), .CP(clk), .CDN(n10), .QN(n55) );
  lanhq1 \hash_I1_reg[14]  ( .E(n20), .D(N255), .Q(hash_I1[14]) );
  dfcrn1 \bits_reg[13]  ( .D(n172), .CP(clk), .CDN(n10), .QN(n56) );
  lanhq1 \hash_I1_reg[13]  ( .E(n21), .D(N254), .Q(hash_I1[13]) );
  dfcrn1 \bits_reg[12]  ( .D(n173), .CP(clk), .CDN(n10), .QN(n57) );
  lanhq1 \hash_I1_reg[12]  ( .E(n21), .D(N253), .Q(hash_I1[12]) );
  dfcrn1 \bits_reg[11]  ( .D(n174), .CP(clk), .CDN(n10), .QN(n58) );
  lanhq1 \hash_I1_reg[11]  ( .E(n21), .D(N252), .Q(hash_I1[11]) );
  dfcrn1 \bits_reg[10]  ( .D(n175), .CP(clk), .CDN(n10), .QN(n59) );
  lanhq1 \hash_I1_reg[10]  ( .E(n21), .D(N251), .Q(hash_I1[10]) );
  dfcrn1 \bits_reg[9]  ( .D(n176), .CP(clk), .CDN(n10), .QN(n60) );
  lanhq1 \hash_I1_reg[9]  ( .E(n21), .D(N250), .Q(hash_I1[9]) );
  dfcrn1 \bits_reg[8]  ( .D(n177), .CP(clk), .CDN(n10), .QN(n61) );
  lanhq1 \hash_I1_reg[8]  ( .E(n21), .D(N249), .Q(hash_I1[8]) );
  dfcrn1 \bits_reg[7]  ( .D(n178), .CP(clk), .CDN(n10), .QN(n62) );
  lanhq1 \hash_I1_reg[7]  ( .E(n21), .D(N248), .Q(hash_I1[7]) );
  dfcrn1 \bits_reg[6]  ( .D(n179), .CP(clk), .CDN(n9), .QN(n63) );
  lanhq1 \hash_I1_reg[6]  ( .E(n21), .D(N247), .Q(hash_I1[6]) );
  dfcrn1 \bits_reg[5]  ( .D(n180), .CP(clk), .CDN(n9), .QN(n64) );
  lanhq1 \hash_I1_reg[5]  ( .E(n21), .D(N246), .Q(hash_I1[5]) );
  dfcrn1 \bits_reg[4]  ( .D(n181), .CP(clk), .CDN(n9), .QN(n65) );
  lanhq1 \hash_I1_reg[4]  ( .E(n22), .D(N245), .Q(hash_I1[4]) );
  dfcrn1 \bits_reg[3]  ( .D(n182), .CP(clk), .CDN(n9), .QN(n66) );
  lanhq1 \hash_I1_reg[3]  ( .E(n22), .D(N244), .Q(hash_I1[3]) );
  dfcrn1 \bits_reg[2]  ( .D(n183), .CP(clk), .CDN(n9), .QN(n67) );
  lanhq1 \hash_I1_reg[2]  ( .E(n22), .D(N243), .Q(hash_I1[2]) );
  dfcrn1 \bits_reg[1]  ( .D(n184), .CP(clk), .CDN(n9), .QN(n68) );
  lanhq1 \hash_I1_reg[1]  ( .E(n22), .D(N242), .Q(hash_I1[1]) );
  dfcrn1 \bits_reg[0]  ( .D(n185), .CP(clk), .CDN(n9), .QN(n69) );
  lanhq1 \hash_I1_reg[0]  ( .E(n22), .D(N241), .Q(hash_I1[0]) );
  an02d1 U68 ( .A1(bit_value), .A2(n102), .Z(n103) );
  an03d1 U69 ( .A1(n223), .A2(n222), .A3(hash_start), .Z(n102) );
  nd04d1 U70 ( .A1(N194), .A2(N193), .A3(n138), .A4(n36), .ZN(n137) );
  an03d1 U73 ( .A1(n141), .A2(n7), .A3(N192), .Z(n138) );
  nr04d1 U75 ( .A1(N159), .A2(n5), .A3(N160), .A4(n146), .ZN(n141) );
  nd04d1 U111 ( .A1(n134), .A2(n224), .A3(n150), .A4(hash_start), .ZN(n148) );
  nr04d1 U114 ( .A1(n100), .A2(hash_A2[5]), .A3(n227), .A4(n153), .ZN(n152) );
  oai22d1 U131 ( .A1(n84), .A2(n85), .B1(n86), .B2(n38), .ZN(n154) );
  oai22d1 U132 ( .A1(n85), .A2(n88), .B1(n89), .B2(n39), .ZN(n155) );
  oai22d1 U133 ( .A1(n85), .A2(n90), .B1(n91), .B2(n40), .ZN(n156) );
  oai22d1 U134 ( .A1(n85), .A2(n92), .B1(n93), .B2(n41), .ZN(n157) );
  oai22d1 U135 ( .A1(n85), .A2(n94), .B1(n95), .B2(n42), .ZN(n158) );
  oai22d1 U136 ( .A1(n85), .A2(n96), .B1(n97), .B2(n43), .ZN(n159) );
  oai22d1 U137 ( .A1(n85), .A2(n98), .B1(n99), .B2(n44), .ZN(n160) );
  oai22d1 U138 ( .A1(n85), .A2(n100), .B1(n101), .B2(n45), .ZN(n161) );
  oai22d1 U139 ( .A1(n84), .A2(n104), .B1(n105), .B2(n46), .ZN(n162) );
  oai22d1 U140 ( .A1(n88), .A2(n104), .B1(n107), .B2(n47), .ZN(n163) );
  oai22d1 U141 ( .A1(n90), .A2(n104), .B1(n108), .B2(n48), .ZN(n164) );
  oai22d1 U142 ( .A1(n92), .A2(n104), .B1(n109), .B2(n49), .ZN(n165) );
  oai22d1 U143 ( .A1(n94), .A2(n104), .B1(n110), .B2(n50), .ZN(n166) );
  oai22d1 U144 ( .A1(n96), .A2(n104), .B1(n111), .B2(n51), .ZN(n167) );
  oai22d1 U145 ( .A1(n98), .A2(n104), .B1(n112), .B2(n52), .ZN(n168) );
  oai22d1 U146 ( .A1(n100), .A2(n104), .B1(n113), .B2(n53), .ZN(n169) );
  oai22d1 U147 ( .A1(n84), .A2(n114), .B1(n115), .B2(n54), .ZN(n170) );
  oai22d1 U148 ( .A1(n88), .A2(n114), .B1(n117), .B2(n55), .ZN(n171) );
  oai22d1 U149 ( .A1(n90), .A2(n114), .B1(n118), .B2(n56), .ZN(n172) );
  oai22d1 U150 ( .A1(n92), .A2(n114), .B1(n119), .B2(n57), .ZN(n173) );
  oai22d1 U151 ( .A1(n94), .A2(n114), .B1(n120), .B2(n58), .ZN(n174) );
  oai22d1 U152 ( .A1(n96), .A2(n114), .B1(n121), .B2(n59), .ZN(n175) );
  oai22d1 U153 ( .A1(n98), .A2(n114), .B1(n122), .B2(n60), .ZN(n176) );
  oai22d1 U154 ( .A1(n100), .A2(n114), .B1(n123), .B2(n61), .ZN(n177) );
  oai22d1 U155 ( .A1(n84), .A2(n124), .B1(n125), .B2(n62), .ZN(n178) );
  oai22d1 U156 ( .A1(n88), .A2(n124), .B1(n127), .B2(n63), .ZN(n179) );
  oai22d1 U157 ( .A1(n90), .A2(n124), .B1(n128), .B2(n64), .ZN(n180) );
  oai22d1 U158 ( .A1(n92), .A2(n124), .B1(n129), .B2(n65), .ZN(n181) );
  oai22d1 U159 ( .A1(n94), .A2(n124), .B1(n130), .B2(n66), .ZN(n182) );
  oai22d1 U160 ( .A1(n96), .A2(n124), .B1(n131), .B2(n67), .ZN(n183) );
  oai22d1 U161 ( .A1(n98), .A2(n124), .B1(n132), .B2(n68), .ZN(n184) );
  oai22d1 U162 ( .A1(n100), .A2(n124), .B1(n133), .B2(n69), .ZN(n185) );
  aon211d1 U163 ( .C1(n135), .C2(n136), .B(n36), .A(n137), .ZN(n186) );
  oai21d1 U164 ( .B1(n135), .B2(n230), .A(n139), .ZN(n187) );
  aoi21d1 U165 ( .B1(n229), .B2(n222), .A(n140), .ZN(n135) );
  aor22d1 U166 ( .A1(n140), .A2(N193), .B1(n229), .B2(n138), .Z(n188) );
  oai21d1 U167 ( .B1(N192), .B2(hash_calc_done), .A(n143), .ZN(n140) );
  oai21d1 U168 ( .B1(n143), .B2(n228), .A(n144), .ZN(n189) );
  aoim21d1 U169 ( .B1(hash_calc_done), .B2(n141), .A(n145), .ZN(n143) );
  or02d0 U170 ( .A1(N162), .A2(N161), .Z(n146) );
  aor22d1 U171 ( .A1(hash_A2[7]), .A2(n145), .B1(N156), .B2(n7), .Z(n190) );
  aor22d1 U172 ( .A1(hash_A2[6]), .A2(n145), .B1(N155), .B2(n7), .Z(n191) );
  aor22d1 U173 ( .A1(hash_A2[5]), .A2(n145), .B1(N154), .B2(n7), .Z(n192) );
  aor22d1 U174 ( .A1(n2), .A2(n145), .B1(N153), .B2(n7), .Z(n193) );
  aor22d1 U175 ( .A1(n4), .A2(n145), .B1(N152), .B2(n7), .Z(n194) );
  aor22d1 U176 ( .A1(hash_A2[2]), .A2(n145), .B1(N151), .B2(n7), .Z(n195) );
  aor22d1 U177 ( .A1(hash_A2[1]), .A2(n145), .B1(N150), .B2(n7), .Z(n196) );
  aor22d1 U178 ( .A1(n6), .A2(n145), .B1(N149), .B2(n7), .Z(n197) );
  aor22d1 U179 ( .A1(hash_A2[8]), .A2(n145), .B1(N157), .B2(n7), .Z(n198) );
  oai21d1 U181 ( .B1(hash_start), .B2(n222), .A(n147), .ZN(n199) );
  oan211d1 U182 ( .C1(N192), .C2(n151), .B(\add_1_root_add_0_root_sub_75/A[3] ), .A(n152), .ZN(n150) );
  or03d0 U183 ( .A1(hash_A2[6]), .A2(hash_A2[8]), .A3(hash_A2[7]), .Z(n153) );
  hash_calc_DW01_inc_1_DW01_inc_4 add_47 ( .A({hash_A2[8:5], n2, n4, 
        hash_A2[2:1], n6}), .SUM({N157, N156, N155, N154, N153, N152, N151, 
        N150, N149}) );
  ah01d1 \add_49/U1_1_1  ( .A(hash_A2[1]), .B(n6), .CO(\add_49/carry[2] ), .S(
        N159) );
  ah01d1 \add_49/U1_1_2  ( .A(hash_A2[2]), .B(\add_49/carry[2] ), .CO(
        \add_49/carry[3] ), .S(N160) );
  ah01d1 \add_49/U1_1_3  ( .A(n4), .B(\add_49/carry[3] ), .CO(
        \add_49/carry[4] ), .S(N161) );
  dfcrq1 \hash_index_reg[2]  ( .D(n187), .CP(clk), .CDN(n9), .Q(N194) );
  dfcrq1 \hash_index_reg[1]  ( .D(n188), .CP(clk), .CDN(n9), .Q(N193) );
  dfcrq1 \hash_index_reg[0]  ( .D(n189), .CP(clk), .CDN(n9), .Q(N192) );
  dfcrq1 hash_calc_done_reg ( .D(n199), .CP(clk), .CDN(n8), .Q(hash_calc_done)
         );
  dfcrq1 \pixel_index_reg[6]  ( .D(n191), .CP(clk), .CDN(n8), .Q(hash_A2[6])
         );
  dfcrq1 \pixel_index_reg[7]  ( .D(n190), .CP(clk), .CDN(n8), .Q(hash_A2[7])
         );
  dfcrq1 \pixel_index_reg[5]  ( .D(n192), .CP(clk), .CDN(n8), .Q(hash_A2[5])
         );
  dfcrq1 \pixel_index_reg[8]  ( .D(n198), .CP(clk), .CDN(n8), .Q(hash_A2[8])
         );
  dfcrq1 \pixel_index_reg[2]  ( .D(n195), .CP(clk), .CDN(n8), .Q(hash_A2[2])
         );
  dfcrq1 \pixel_index_reg[1]  ( .D(n196), .CP(clk), .CDN(n8), .Q(hash_A2[1])
         );
  dfcrq1 \pixel_index_reg[4]  ( .D(n193), .CP(clk), .CDN(n8), .Q(hash_A2[4])
         );
  dfcrq1 \pixel_index_reg[3]  ( .D(n194), .CP(clk), .CDN(n8), .Q(hash_A2[3])
         );
  dfcrq1 \pixel_index_reg[0]  ( .D(n197), .CP(clk), .CDN(n8), .Q(hash_A2[0])
         );
  inv0d0 U7 ( .I(hash_A2[0]), .ZN(n5) );
  inv0d0 U8 ( .I(hash_A2[3]), .ZN(n3) );
  inv0d0 U9 ( .I(hash_A2[4]), .ZN(n1) );
  buffd1 U19 ( .I(n23), .Z(n21) );
  buffd1 U20 ( .I(n23), .Z(n20) );
  buffd1 U21 ( .I(n23), .Z(n22) );
  buffd1 U22 ( .I(n37), .Z(n19) );
  buffd1 U23 ( .I(N228), .Z(n37) );
  buffd1 U24 ( .I(N228), .Z(n23) );
  nd03d1 U25 ( .A1(n4), .A2(n102), .A3(n2), .ZN(n87) );
  nd03d1 U26 ( .A1(n102), .A2(n1), .A3(n4), .ZN(n116) );
  nd03d1 U27 ( .A1(n102), .A2(n3), .A3(n2), .ZN(n106) );
  nd02d1 U28 ( .A1(n134), .A2(n102), .ZN(n126) );
  nr02d1 U29 ( .A1(n4), .A2(n2), .ZN(n134) );
  nd02d1 U30 ( .A1(n149), .A2(n148), .ZN(N228) );
  inv0d0 U31 ( .I(n16), .ZN(n14) );
  inv0d0 U32 ( .I(n17), .ZN(n13) );
  nd03d1 U33 ( .A1(n4), .A2(n1), .A3(n103), .ZN(n114) );
  nd03d1 U34 ( .A1(n2), .A2(n3), .A3(n103), .ZN(n104) );
  nd03d1 U35 ( .A1(n2), .A2(n4), .A3(n103), .ZN(n85) );
  nd02d1 U36 ( .A1(n134), .A2(n103), .ZN(n124) );
  inv0d0 U37 ( .I(n1), .ZN(n2) );
  inv0d0 U38 ( .I(n3), .ZN(n4) );
  inv0d0 U39 ( .I(n5), .ZN(n6) );
  nd03d1 U40 ( .A1(n225), .A2(n226), .A3(n5), .ZN(n100) );
  nd03d1 U41 ( .A1(n225), .A2(n226), .A3(n6), .ZN(n98) );
  nd02d1 U42 ( .A1(n152), .A2(hash_start), .ZN(n149) );
  buffd1 U43 ( .I(n231), .Z(n8) );
  buffd1 U44 ( .I(n231), .Z(n9) );
  buffd1 U45 ( .I(n231), .Z(n10) );
  buffd1 U46 ( .I(n231), .Z(n11) );
  buffd1 U47 ( .I(n18), .Z(n15) );
  buffd1 U48 ( .I(n18), .Z(n16) );
  buffd1 U49 ( .I(n18), .Z(n17) );
  inv0d0 U50 ( .I(n83), .ZN(n220) );
  buffd1 U51 ( .I(n231), .Z(n12) );
  nd02d1 U52 ( .A1(n229), .A2(n230), .ZN(n151) );
  nd02d1 U53 ( .A1(n222), .A2(n230), .ZN(n136) );
  nd03d1 U54 ( .A1(n138), .A2(n230), .A3(N193), .ZN(n139) );
  nd03d1 U55 ( .A1(n7), .A2(n228), .A3(n141), .ZN(n144) );
  inv0d0 U56 ( .I(N192), .ZN(n228) );
  nr02d1 U57 ( .A1(n100), .A2(n116), .ZN(n123) );
  nr02d1 U58 ( .A1(n100), .A2(n106), .ZN(n113) );
  nr02d1 U59 ( .A1(n98), .A2(n116), .ZN(n122) );
  nr02d1 U60 ( .A1(n96), .A2(n116), .ZN(n121) );
  nr02d1 U61 ( .A1(n94), .A2(n116), .ZN(n120) );
  nr02d1 U62 ( .A1(n92), .A2(n116), .ZN(n119) );
  nr02d1 U63 ( .A1(n90), .A2(n116), .ZN(n118) );
  nr02d1 U64 ( .A1(n88), .A2(n116), .ZN(n117) );
  nr02d1 U65 ( .A1(n84), .A2(n116), .ZN(n115) );
  nr02d1 U66 ( .A1(n98), .A2(n106), .ZN(n112) );
  nr02d1 U67 ( .A1(n96), .A2(n106), .ZN(n111) );
  nr02d1 U71 ( .A1(n94), .A2(n106), .ZN(n110) );
  nr02d1 U72 ( .A1(n92), .A2(n106), .ZN(n109) );
  nr02d1 U74 ( .A1(n90), .A2(n106), .ZN(n108) );
  nr02d1 U76 ( .A1(n88), .A2(n106), .ZN(n107) );
  nr02d1 U77 ( .A1(n84), .A2(n106), .ZN(n105) );
  oai21d1 U78 ( .B1(hash_calc_done), .B2(n223), .A(hash_start), .ZN(n145) );
  buffd1 U79 ( .I(n142), .Z(n7) );
  nr02d1 U80 ( .A1(n145), .A2(hash_calc_done), .ZN(n142) );
  nr02d1 U81 ( .A1(n87), .A2(n84), .ZN(n86) );
  nr02d1 U82 ( .A1(n87), .A2(n100), .ZN(n101) );
  nr02d1 U83 ( .A1(n87), .A2(n98), .ZN(n99) );
  nr02d1 U84 ( .A1(n87), .A2(n96), .ZN(n97) );
  nr02d1 U85 ( .A1(n87), .A2(n94), .ZN(n95) );
  nr02d1 U86 ( .A1(n87), .A2(n92), .ZN(n93) );
  nr02d1 U87 ( .A1(n87), .A2(n90), .ZN(n91) );
  nr02d1 U88 ( .A1(n87), .A2(n88), .ZN(n89) );
  nr02d1 U89 ( .A1(n100), .A2(n126), .ZN(n133) );
  nr02d1 U90 ( .A1(n98), .A2(n126), .ZN(n132) );
  nr02d1 U91 ( .A1(n96), .A2(n126), .ZN(n131) );
  nr02d1 U92 ( .A1(n94), .A2(n126), .ZN(n130) );
  nr02d1 U93 ( .A1(n92), .A2(n126), .ZN(n129) );
  nr02d1 U94 ( .A1(n90), .A2(n126), .ZN(n128) );
  nr02d1 U95 ( .A1(n88), .A2(n126), .ZN(n127) );
  nr02d1 U96 ( .A1(n84), .A2(n126), .ZN(n125) );
  inv0d0 U97 ( .I(hash_calc_done), .ZN(n222) );
  inv0d0 U98 ( .I(hash_A2[8]), .ZN(n223) );
  nd03d1 U99 ( .A1(hash_start), .A2(n222), .A3(hash_A2[8]), .ZN(n147) );
  inv0d0 U100 ( .I(hash_A2[1]), .ZN(n225) );
  inv0d0 U101 ( .I(hash_A2[2]), .ZN(n226) );
  nd03d1 U102 ( .A1(n5), .A2(n226), .A3(hash_A2[1]), .ZN(n96) );
  nd03d1 U103 ( .A1(n5), .A2(n225), .A3(hash_A2[2]), .ZN(n92) );
  nd03d1 U104 ( .A1(hash_A2[1]), .A2(n5), .A3(hash_A2[2]), .ZN(n88) );
  nd03d1 U105 ( .A1(n6), .A2(n225), .A3(hash_A2[2]), .ZN(n90) );
  nd03d1 U106 ( .A1(n6), .A2(n226), .A3(hash_A2[1]), .ZN(n94) );
  nd03d1 U107 ( .A1(hash_A2[1]), .A2(n6), .A3(hash_A2[2]), .ZN(n84) );
  inv0d0 U108 ( .I(N193), .ZN(n229) );
  inv0d0 U109 ( .I(N194), .ZN(n230) );
  inv0d0 U110 ( .I(n134), .ZN(n227) );
  inv0d0 U112 ( .I(n75), .ZN(n216) );
  inv0d0 U113 ( .I(hash_O2[0]), .ZN(n211) );
  inv0d0 U115 ( .I(reset), .ZN(n231) );
  inv0d0 U116 ( .I(n148), .ZN(n18) );
  inv0d0 U117 ( .I(n100), .ZN(n224) );
  inv0d0 U118 ( .I(n80), .ZN(n221) );
  nr02d1 U119 ( .A1(n69), .A2(n148), .ZN(N241) );
  nr02d1 U120 ( .A1(n68), .A2(n148), .ZN(N242) );
  nr02d1 U121 ( .A1(n67), .A2(n14), .ZN(N243) );
  nr02d1 U122 ( .A1(n66), .A2(n14), .ZN(N244) );
  nr02d1 U123 ( .A1(n65), .A2(n14), .ZN(N245) );
  nr02d1 U124 ( .A1(n64), .A2(n14), .ZN(N246) );
  nr02d1 U125 ( .A1(n63), .A2(n14), .ZN(N247) );
  nr02d1 U126 ( .A1(n62), .A2(n14), .ZN(N248) );
  nr02d1 U127 ( .A1(n61), .A2(n14), .ZN(N249) );
  nr02d1 U128 ( .A1(n60), .A2(n14), .ZN(N250) );
  nr02d1 U129 ( .A1(n59), .A2(n14), .ZN(N251) );
  nr02d1 U130 ( .A1(n58), .A2(n14), .ZN(N252) );
  nr02d1 U180 ( .A1(n57), .A2(n13), .ZN(N253) );
  nr02d1 U184 ( .A1(n56), .A2(n13), .ZN(N254) );
  nr02d1 U185 ( .A1(n55), .A2(n13), .ZN(N255) );
  nr02d1 U186 ( .A1(n54), .A2(n13), .ZN(N256) );
  nr02d1 U187 ( .A1(n53), .A2(n13), .ZN(N257) );
  nr02d1 U188 ( .A1(n52), .A2(n13), .ZN(N258) );
  nr02d1 U189 ( .A1(n51), .A2(n13), .ZN(N259) );
  nr02d1 U190 ( .A1(n50), .A2(n13), .ZN(N260) );
  nr02d1 U191 ( .A1(n49), .A2(n13), .ZN(N261) );
  nr02d1 U192 ( .A1(n48), .A2(n13), .ZN(N262) );
  nr02d1 U193 ( .A1(n47), .A2(n148), .ZN(N263) );
  nr02d1 U194 ( .A1(n46), .A2(n148), .ZN(N264) );
  nr02d1 U195 ( .A1(n45), .A2(n148), .ZN(N265) );
  nr02d1 U196 ( .A1(n44), .A2(n148), .ZN(N266) );
  nr02d1 U197 ( .A1(n43), .A2(n148), .ZN(N267) );
  nr02d1 U198 ( .A1(n42), .A2(n148), .ZN(N268) );
  nr02d1 U199 ( .A1(n41), .A2(n148), .ZN(N269) );
  nr02d1 U200 ( .A1(n40), .A2(n148), .ZN(N270) );
  nr02d1 U201 ( .A1(n39), .A2(n148), .ZN(N271) );
  nr02d1 U202 ( .A1(n38), .A2(n148), .ZN(N272) );
  inv0d0 U203 ( .I(n36), .ZN(\add_1_root_add_0_root_sub_75/A[3] ) );
  inv0d0 U204 ( .I(sum[12]), .ZN(n217) );
  inv0d0 U205 ( .I(hash_O2[3]), .ZN(n213) );
  inv0d0 U206 ( .I(sum[9]), .ZN(n215) );
  inv0d0 U207 ( .I(hash_O2[7]), .ZN(n214) );
  inv0d0 U208 ( .I(sum[13]), .ZN(n218) );
  inv0d0 U209 ( .I(hash_O2[2]), .ZN(n212) );
  inv0d0 U210 ( .I(sum[14]), .ZN(n219) );
  xr02d1 U211 ( .A1(N203), .A2(\add_0_root_add_0_root_sub_75/carry[11] ), .Z(
        N227) );
  an02d0 U212 ( .A1(\add_0_root_add_0_root_sub_75/carry[10] ), .A2(N202), .Z(
        \add_0_root_add_0_root_sub_75/carry[11] ) );
  xr02d1 U213 ( .A1(N202), .A2(\add_0_root_add_0_root_sub_75/carry[10] ), .Z(
        N226) );
  an02d0 U214 ( .A1(\add_0_root_add_0_root_sub_75/carry[9] ), .A2(N201), .Z(
        \add_0_root_add_0_root_sub_75/carry[10] ) );
  xr02d1 U215 ( .A1(N201), .A2(\add_0_root_add_0_root_sub_75/carry[9] ), .Z(
        N225) );
  an02d0 U216 ( .A1(\add_0_root_add_0_root_sub_75/carry[8] ), .A2(N200), .Z(
        \add_0_root_add_0_root_sub_75/carry[9] ) );
  xr02d1 U217 ( .A1(N200), .A2(\add_0_root_add_0_root_sub_75/carry[8] ), .Z(
        N224) );
  or02d0 U218 ( .A1(N199), .A2(\add_0_root_add_0_root_sub_75/carry[7] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[8] ) );
  xn02d1 U219 ( .A1(\add_0_root_add_0_root_sub_75/carry[7] ), .A2(N199), .ZN(
        N223) );
  or02d0 U220 ( .A1(N198), .A2(\add_0_root_add_0_root_sub_75/carry[6] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[7] ) );
  xn02d1 U221 ( .A1(\add_0_root_add_0_root_sub_75/carry[6] ), .A2(N198), .ZN(
        N222) );
  or02d0 U222 ( .A1(N197), .A2(\add_0_root_add_0_root_sub_75/carry[5] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[6] ) );
  xn02d1 U223 ( .A1(\add_0_root_add_0_root_sub_75/carry[5] ), .A2(N197), .ZN(
        N221) );
  or02d0 U224 ( .A1(N196), .A2(\add_0_root_add_0_root_sub_75/carry[4] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[5] ) );
  xn02d1 U225 ( .A1(\add_0_root_add_0_root_sub_75/carry[4] ), .A2(N196), .ZN(
        N220) );
  or02d0 U226 ( .A1(N195), .A2(\add_0_root_add_0_root_sub_75/carry[3] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[4] ) );
  xn02d1 U227 ( .A1(\add_0_root_add_0_root_sub_75/carry[3] ), .A2(N195), .ZN(
        N219) );
  or02d0 U228 ( .A1(N194), .A2(\add_0_root_add_0_root_sub_75/carry[2] ), .Z(
        \add_0_root_add_0_root_sub_75/carry[3] ) );
  xn02d1 U229 ( .A1(\add_0_root_add_0_root_sub_75/carry[2] ), .A2(N194), .ZN(
        N218) );
  or02d0 U230 ( .A1(N193), .A2(N192), .Z(
        \add_0_root_add_0_root_sub_75/carry[2] ) );
  xn02d1 U231 ( .A1(N192), .A2(N193), .ZN(N217) );
  xr02d1 U232 ( .A1(image_header[8]), .A2(
        \add_1_root_add_0_root_sub_75/carry[11] ), .Z(N203) );
  an02d0 U233 ( .A1(\add_1_root_add_0_root_sub_75/carry[10] ), .A2(
        image_header[7]), .Z(\add_1_root_add_0_root_sub_75/carry[11] ) );
  xr02d1 U234 ( .A1(image_header[7]), .A2(
        \add_1_root_add_0_root_sub_75/carry[10] ), .Z(N202) );
  an02d0 U235 ( .A1(\add_1_root_add_0_root_sub_75/carry[9] ), .A2(
        image_header[6]), .Z(\add_1_root_add_0_root_sub_75/carry[10] ) );
  xr02d1 U236 ( .A1(image_header[6]), .A2(
        \add_1_root_add_0_root_sub_75/carry[9] ), .Z(N201) );
  an02d0 U237 ( .A1(\add_1_root_add_0_root_sub_75/carry[8] ), .A2(
        image_header[5]), .Z(\add_1_root_add_0_root_sub_75/carry[9] ) );
  xr02d1 U238 ( .A1(image_header[5]), .A2(
        \add_1_root_add_0_root_sub_75/carry[8] ), .Z(N200) );
  an02d0 U239 ( .A1(\add_1_root_add_0_root_sub_75/carry[7] ), .A2(
        image_header[4]), .Z(\add_1_root_add_0_root_sub_75/carry[8] ) );
  xr02d1 U240 ( .A1(image_header[4]), .A2(
        \add_1_root_add_0_root_sub_75/carry[7] ), .Z(N199) );
  an02d0 U241 ( .A1(\add_1_root_add_0_root_sub_75/carry[6] ), .A2(
        image_header[3]), .Z(\add_1_root_add_0_root_sub_75/carry[7] ) );
  xr02d1 U242 ( .A1(image_header[3]), .A2(
        \add_1_root_add_0_root_sub_75/carry[6] ), .Z(N198) );
  an02d0 U243 ( .A1(\add_1_root_add_0_root_sub_75/carry[5] ), .A2(
        image_header[2]), .Z(\add_1_root_add_0_root_sub_75/carry[6] ) );
  xr02d1 U244 ( .A1(image_header[2]), .A2(
        \add_1_root_add_0_root_sub_75/carry[5] ), .Z(N197) );
  an02d0 U245 ( .A1(\add_1_root_add_0_root_sub_75/carry[4] ), .A2(
        image_header[1]), .Z(\add_1_root_add_0_root_sub_75/carry[5] ) );
  xr02d1 U246 ( .A1(image_header[1]), .A2(
        \add_1_root_add_0_root_sub_75/carry[4] ), .Z(N196) );
  an02d0 U247 ( .A1(\add_1_root_add_0_root_sub_75/A[3] ), .A2(image_header[0]), 
        .Z(\add_1_root_add_0_root_sub_75/carry[4] ) );
  xr02d1 U248 ( .A1(image_header[0]), .A2(\add_1_root_add_0_root_sub_75/A[3] ), 
        .Z(N195) );
  xr02d1 U249 ( .A1(\add_49/carry[4] ), .A2(n2), .Z(N162) );
  nr04d0 U250 ( .A1(n4), .A2(hash_A2[2]), .A3(hash_A2[1]), .A4(n6), .ZN(n71)
         );
  nr04d0 U251 ( .A1(hash_A2[7]), .A2(hash_A2[6]), .A3(hash_A2[5]), .A4(n2), 
        .ZN(n70) );
  oaim21d1 U252 ( .B1(n71), .B2(n70), .A(hash_A2[8]), .ZN(N273) );
  nr03d0 U253 ( .A1(hash_O2[14]), .A2(hash_O2[16]), .A3(hash_O2[15]), .ZN(n210) );
  nr04d0 U254 ( .A1(hash_O2[20]), .A2(hash_O2[19]), .A3(hash_O2[18]), .A4(
        hash_O2[17]), .ZN(n209) );
  or02d0 U255 ( .A1(hash_O2[5]), .A2(n218), .Z(n79) );
  an02d0 U256 ( .A1(sum[11]), .A2(n213), .Z(n73) );
  nr03d0 U257 ( .A1(n73), .A2(sum[10]), .A3(n212), .ZN(n72) );
  aoim21d1 U258 ( .B1(sum[11]), .B2(n213), .A(n72), .ZN(n75) );
  aon211d1 U259 ( .C1(sum[10]), .C2(n212), .B(n73), .A(n75), .ZN(n74) );
  oai211d1 U260 ( .C1(hash_O2[4]), .C2(n217), .A(n79), .B(n74), .ZN(n201) );
  aoim22d1 U261 ( .A1(sum[8]), .A2(n211), .B1(n215), .B2(hash_O2[1]), .Z(n76)
         );
  aoi211d1 U262 ( .C1(hash_O2[1]), .C2(n215), .A(n216), .B(n76), .ZN(n200) );
  nd02d0 U263 ( .A1(sum[15]), .A2(n214), .ZN(n77) );
  oai21d1 U264 ( .B1(hash_O2[6]), .B2(n219), .A(n77), .ZN(n83) );
  nd03d0 U265 ( .A1(n77), .A2(n219), .A3(hash_O2[6]), .ZN(n78) );
  oai21d1 U266 ( .B1(sum[15]), .B2(n214), .A(n78), .ZN(n81) );
  aoi321d1 U267 ( .C1(hash_O2[4]), .C2(n217), .C3(n79), .B1(n218), .B2(
        hash_O2[5]), .A(n81), .ZN(n80) );
  oan211d1 U268 ( .C1(n220), .C2(n81), .B(n221), .A(hash_O2[10]), .ZN(n82) );
  oai31d1 U269 ( .B1(n201), .B2(n200), .B3(n83), .A(n82), .ZN(n202) );
  nr04d0 U270 ( .A1(n202), .A2(hash_O2[11]), .A3(hash_O2[13]), .A4(hash_O2[12]), .ZN(n208) );
  nr03d0 U271 ( .A1(hash_O2[21]), .A2(hash_O2[23]), .A3(hash_O2[22]), .ZN(n206) );
  nr03d0 U272 ( .A1(hash_O2[24]), .A2(hash_O2[26]), .A3(hash_O2[25]), .ZN(n205) );
  nr03d0 U273 ( .A1(hash_O2[27]), .A2(hash_O2[29]), .A3(hash_O2[28]), .ZN(n204) );
  nr04d0 U274 ( .A1(hash_O2[9]), .A2(hash_O2[8]), .A3(hash_O2[31]), .A4(
        hash_O2[30]), .ZN(n203) );
  an04d0 U275 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .Z(n207) );
  nd04d0 U276 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(N274) );
endmodule


module reordering_DW01_inc_0_DW01_inc_2 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ah01d1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ah01d1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ah01d1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ah01d1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ah01d1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ah01d1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ah01d1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  inv0d0 U1 ( .I(A[0]), .ZN(SUM[0]) );
  xr02d1 U2 ( .A1(carry[8]), .A2(A[8]), .Z(SUM[8]) );
endmodule


module reordering_DW01_add_9 ( A, B, CI, SUM, CO );
  input [8:0] A;
  input [8:0] B;
  output [8:0] SUM;
  input CI;
  output CO;
  wire   n2;
  wire   [8:1] carry;

  ad01d0 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  ad01d0 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  ad01d0 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  ad01d0 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  ad01d0 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  ad01d0 U1_1 ( .A(A[1]), .B(B[1]), .CI(n2), .CO(carry[2]), .S(SUM[1]) );
  an02d1 U1 ( .A1(B[7]), .A2(carry[7]), .Z(SUM[8]) );
  an02d1 U2 ( .A1(B[0]), .A2(A[0]), .Z(n2) );
  xr02d1 U3 ( .A1(B[0]), .A2(A[0]), .Z(SUM[0]) );
  xr02d1 U4 ( .A1(B[7]), .A2(carry[7]), .Z(SUM[7]) );
endmodule


module reordering_DW01_inc_1_DW01_inc_6 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ah01d1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ah01d1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ah01d1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ah01d1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ah01d1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ah01d1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ah01d1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  inv0d0 U1 ( .I(A[0]), .ZN(SUM[0]) );
  xr02d1 U2 ( .A1(carry[8]), .A2(A[8]), .Z(SUM[8]) );
endmodule


module reordering ( clk, reset, num_images, reorder_start, temp_new_reference, 
        new_reference_is_done, count_image, last_image, finish_reordering, 
        reorder_O1, reorder_O2, reorder_A1, reorder_A2, reorder_WEB1, 
        reorder_WEB2 );
  input [8:0] num_images;
  output [8:0] temp_new_reference;
  output [8:0] count_image;
  output [8:0] last_image;
  input [31:0] reorder_O1;
  input [31:0] reorder_O2;
  output [11:0] reorder_A1;
  output [11:0] reorder_A2;
  input clk, reset, reorder_start;
  output new_reference_is_done, finish_reordering, reorder_WEB1, reorder_WEB2;
  wire   N3179, N3180, N3181, N3182, reading_current, reading_compare,
         hashes_ready, compare_in_progress, distance_ready, finish_flag, N3187,
         N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3231,
         N3232, N3233, N3234, N3235, N3237, N3238, N3239, N3843, N3844, N3845,
         N3846, N3847, N3848, N3849, N3850, N3851, N3877, N3878, N3879, N3880,
         N3881, N3882, N3883, N3884, N3885, N3886, N3887, N3914, N3915, N3972,
         N3973, N3974, N3975, N3976, N3978, N3979, N3980, N4002, N4003, N4004,
         N4010, N4011, N4012, N4013, N4652, N4653, N4654, N4655, N4656, N4657,
         N4658, N4659, N4660, N4688, N4689, N4690, N4691, N4692, N4693, N4694,
         N4695, N4696, N4723, N4724, N4760, N4764, N4765, N4766, N4767, N4768,
         N4769, N4770, N4771, N4772, N4773, N4774, N4775, N4776, N4777, N4778,
         N4779, N4780, N4781, N4782, N4783, N4784, N4785, N4786, N4787, N4788,
         N4789, N4790, N4791, N4792, N4793, N4794, N4795, N4796, N4797, N4798,
         N4799, N4800, N4801, N4802, N4803, N4804, N4805, N4806, N4807, N4808,
         N4809, N4810, N4811, N4812, N4813, N4814, N4815, N4816, N4817, N4818,
         N4819, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828,
         N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838,
         N4839, N4840, N4841, N4842, N4843, N4844, N4845, N4846, N4847, N4848,
         N4849, N4850, N4851, N4852, N4853, N4854, N4855, N4856, N4857, N4858,
         N4859, N4860, N4861, N4862, N4863, N4864, N4865, N4866, N4867, N4868,
         N4869, N4870, N4871, N4872, N4873, N4874, N4875, N4876, N4877, N4878,
         N4879, N4880, N4881, N4882, N4883, N4884, N4885, N4886, N4887, N4888,
         N4889, N4890, N4891, N4892, N4893, N4894, N4895, N4896, N4897, N4898,
         N4899, N4900, N4901, N4902, N4903, N4904, N4905, N4906, N4907, N4908,
         N4909, N4910, N4911, N4912, N4913, N4914, N4915, N4916, N4917, N4918,
         N4919, N4920, N4921, N4922, N4923, N4924, N4925, N4926, N4927, N4928,
         N4929, N4930, N4931, N4932, N4933, N4934, N4935, N4936, N4937, N4938,
         N4939, N4940, N4941, N4942, N4943, N4944, N4945, N4946, N4947, N4948,
         N4949, N4950, N4951, N4952, N4953, N4954, N4955, N4956, N4957, N4958,
         N4959, N4960, N4961, N4962, N4963, N4964, N4965, N4966, N4967, N4968,
         N4969, N4970, N4971, N4972, N4973, N4974, N4975, N4976, N4977, N4978,
         N4979, N4980, N4981, N4982, N4983, N4984, N4985, N4986, N4987, N4988,
         N4989, N4990, N4991, N4992, N4993, N4994, N4995, N4996, N4997, N4998,
         N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008,
         N5009, N5010, N5011, N5012, N5013, N5014, N5015, N5016, N5017, N5018,
         N5019, N5020, N5021, N5022, N5023, N5024, N5025, N5026, N5027, N5028,
         N5029, N5070, N5071, N5072, N5073, N5074, N5076, N5077, N5078, N5108,
         N5109, N5110, N5111, N5113, N5114, N5115, N5116, N5117, N5118, N5119,
         N5120, N5121, N5122, N5285, N6837, N6838, N6839, N6840, N6841, N6842,
         N6843, N6844, N6845, N6867, N6869, N6870, N6871, N6872, N6873, N6874,
         N6875, N7997, N8001, N8008, N8016, N8025, N8034, N8044, N8054, N8064,
         N8074, N8085, N8096, N8107, N8129, N8151, N8162, N8174, N8186, N8198,
         N8210, N8234, N8246, N8258, N8270, N8282, N8294, N8306, N8318, N8330,
         N8342, N8354, N8367, N8380, N8393, N8406, N8432, N8445, N8458, N8471,
         N8484, N8497, N8510, N8523, N8536, N8549, N8562, N8575, N8601, N8614,
         N8627, N8640, N8653, N8666, N8679, N8692, N8705, N8718, N8731, N8744,
         N8770, N8784, N8798, N8812, N8826, N8840, N8854, N8868, N8882, N8896,
         N8910, N8924, N8938, N8952, N8980, N8994, N9008, N9022, N9036, N9050,
         N9064, N9078, N9092, N9106, N9120, N9134, N9148, N9162, N9176, N9190,
         N9204, N9218, N9232, N9246, N9260, N9274, N9288, N9302, N9316, N9330,
         N9344, N9358, N9372, N9386, N9400, N9414, N9428, N9442, N9456, N9470,
         N9484, N9498, N9512, N9526, N9540, N9554, N9568, N9582, N9596, N9610,
         N9624, N9638, N9652, N9666, N9681, N9696, N9711, N9726, N9741, N9756,
         N9786, N9801, N9816, N9831, N9846, N9861, N9876, N9891, N9906, N9921,
         N9936, N9951, N9966, N9981, N9996, N10011, N10026, N10041, N10056,
         N10071, N10086, N10101, N10131, N10146, N10161, N10176, N10191,
         N10206, N10221, N10236, N10251, N10266, N10281, N10296, N10311,
         N10326, N10341, N10371, N10386, N10401, N10416, N10431, N10446,
         N10461, N10476, N10491, N10506, N10521, N10536, N10551, N10566,
         N10581, N10596, N10611, N10626, N10641, N10656, N10671, N10686,
         N10701, N10716, N10731, N10746, N10761, N10776, N10791, N10806,
         N10821, N10836, N10851, N10866, N10881, N10896, N10911, N10926,
         N10941, N10956, N10971, N10986, N11001, N11016, N11031, N11046,
         N11061, N11076, N11091, N11106, N11121, N11136, N11151, N11166,
         N11181, N11196, N11211, N11226, N11241, N11256, N11271, N11286,
         N11301, N11316, N11331, N11346, N11376, N11391, N11406, N11421,
         N11436, N11451, N11466, N11481, N11496, N11511, N11526, N11541,
         N11556, N11571, N11586, N11602, N11618, N11634, N11650, N11666,
         N11682, N11698, N11714, N11730, N11746, N11762, N11778, N11794,
         N11810, N11826, N11842, N11858, N11874, N11890, N11906, N11922,
         N11938, N11954, N11970, N11986, N12002, N12018, N12034, N12050,
         N12066, N12082, N12098, N12114, N12130, N12146, N12162, N12178,
         N12194, N12210, N12226, N12242, N12258, N12274, N12290, N12306,
         N12322, N12338, N12354, N12370, N12386, N12402, N12418, N12434,
         N12450, N12466, N12482, N12498, N12514, N12530, N12546, N12562,
         N12594, N12610, N12626, N12658, N12674, N12690, N12706, N12722,
         N12738, N12754, N12786, N12802, N12818, N12850, N12866, N12882,
         N12898, N12914, N12930, N12946, N12962, N12978, N12994, N13010,
         N13026, N13042, N13058, N13074, N13090, N13106, N13122, N13138,
         N13170, N13186, N13202, N13234, N13250, N13266, N13282, N13298,
         N13314, N13330, N13346, N13362, N13378, N13394, N13410, N13426,
         N13442, N13458, N13490, N13506, N13522, N13538, N13554, N13570,
         N13586, N13602, N13650, N13666, N13682, N13714, N13730, N13746,
         N13762, N13778, N13794, N13810, N13826, N13858, N13874, N13890,
         N13906, N13922, N13938, N13954, N13970, N13986, N14002, N14018,
         N14034, N14050, N14066, N14082, N14098, N14114, N14130, N14146,
         N14162, N14178, N14194, N14210, N14226, N14242, N14258, N14274,
         N14290, N14306, N14322, N14338, N14354, N14370, N14386, N14402,
         N14418, N14434, N14450, N14466, N14482, N14498, N14514, N14530,
         N14546, N14562, N14578, N14594, N14610, N14626, N14658, N14690,
         N14706, N14722, N14738, N14754, N14770, N14802, N14834, N14850,
         N14866, N14882, N14930, N14946, N14962, N14994, N15010, N15026,
         N15042, N15058, N15074, N15090, N15106, N15122, N15154, N15170,
         N15186, N15202, N15218, N15234, N15250, N15266, N15282, N15298,
         N15314, N15330, N15346, N15362, N15378, N15394, N15410, N15442,
         N15458, N15474, N15490, N15522, N15538, N15554, N15570, N15586,
         N15602, N15618, N15633, N26357, N26358, N26359, N26360, N26361,
         N26362, N26363, N26364, N26365, N26366, N26480, N26489, n3578, n3579,
         n3580, n3581, n3583, n3584, n3585, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3620, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3651, n3652, n3654, n3655, n3656, n3657,
         n3658, n3661, n3662, n3663, n3666, n3667, n3669, n3670, n3671, n3673,
         n3674, n3676, n3677, n3680, n3682, n3683, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3693, n3694, n3695, n3696, n3697, n3698, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3709, n3710, n3711, n3713,
         n3714, n3716, n3718, n3720, n3722, n3724, n3726, n3727, n3729, n3731,
         n3733, n3735, n3737, n3739, n3741, n3743, n3745, n3747, n3749, n3750,
         n3752, n3754, n3756, n3758, n3760, n3762, n3763, n3765, n3767, n3768,
         n3794, n3796, n3797, n3825, n3827, n3855, n3884, n3885, n3918, n3948,
         n3949, n3980, n4010, n4011, n4040, n4069, n4100, n4131, n4162, n4192,
         n4193, n4194, n4197, n4198, n4200, n4202, n4204, n4206, n4208, n4211,
         n4212, n4221, n4234, n4235, n4236, n4237, n4240, n4241, n4242, n4245,
         n4254, n4258, n4327, n4329, n4332, n4335, n4336, n4337, n4340, n4343,
         n4344, n4345, n4349, n4350, n4353, n4354, n4355, n4356, n4358, n4359,
         n4360, n4362, n4363, n4364, n4367, n4370, n4371, n4372, n4375, n4377,
         n4378, n4379, n4380, n4381, n4382, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4394, n4395, n4398, n4399, n4400, n4401, n4402, n4403,
         n4407, n4409, n4410, n4412, n4413, n4414, n4415, n4417, n4418, n4420,
         n4422, n4424, n4425, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4440, n4442, n4443, n4445, n4446, n4447, n4448, n4449, n4452,
         n4453, n4454, n4455, n4456, n4458, n4460, n4461, n4463, n4465, n4466,
         n4467, n4468, n4469, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4492, n4494, n4495, n4496, n4498, n4499, n4500, n4501, n4502,
         n4504, n4505, n4507, n4508, n4509, n4511, n4513, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4525, n4526, n4527, n4528, n4529,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4550, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4562, n4563, n4564,
         n4565, n4566, n4567, n4569, n4570, n4571, n4573, n4574, n4577, n4578,
         n4579, n4581, n4582, n4583, n4584, n4585, n4586, n4588, n4589, n4591,
         n4592, n4593, n4594, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4605, n4606, n4607, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4629, n4630, n4631, n4632, n4634, n4636, n4637, n4638,
         n4639, n4641, n4642, n4643, n4644, n4645, n4647, n4648, n4650, n4651,
         n4652, n4654, n4655, n4657, n4658, n4659, n4660, n4661, n4662, n4664,
         n4665, n4666, n4667, n4669, n4670, n4671, n4672, n4673, n4674, n4676,
         n4678, n4679, n4680, n4682, n4684, n4685, n4686, n4687, n4688, n4690,
         n4694, n4695, n4696, n4697, n4699, n4700, n4701, n4702, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4712, n4713, n4714, n4715, n4716,
         n4717, n4718, n4720, n4721, n4722, n4723, n4724, n4726, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4736, n4737, n4738, n4739, n4740,
         n4741, n4743, n4744, n4748, n4749, n4750, n4752, n4753, n4755, n4756,
         n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4768,
         n4769, n4770, n4772, n4773, n4774, n4775, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4790, n4791,
         n4792, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4817, n4818, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4828, n4829, n4830, n4831, n4833, n4834, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4845, n4846, n4848, n4849,
         n4850, n4851, n4852, n4853, n4855, n4856, n4857, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4867, n4868, n4869, n4870, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4882, n4883, n4884,
         n4885, n4887, n4888, n4891, n4892, n4893, n4896, n4897, n4898, n4899,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4914, n4916, n4917, n4918, n4919, n4920, n4921, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4940, n4942, n4943, n4945, n4947, n4950, n4952,
         n4953, n4955, n4956, n4960, n4961, n4963, n4964, n4967, n4968, n4969,
         n4970, n4971, n4972, n4975, n4977, n4978, n4979, n4981, n4982, n4983,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n5000, n5001, n5002, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5045, n5047, n5048, n5050, n5051, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5062, n5064, n5065, n5066, n5067,
         n5069, n5070, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5094, n5095, n5097, n5099, n5100, n5102, n5103, n5105,
         n5107, n5108, n5109, n5111, n5112, n5114, n5115, n5116, n5117, n5119,
         n5120, n5121, n5122, n5123, n5125, n5127, n5128, n5130, n5131, n5132,
         n5133, n5134, n5135, n5137, n5138, n5139, n5141, n5143, n5144, n5147,
         n5148, n5149, n5150, n5151, n5153, n5154, n5155, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5166, n5167, n5169, n5170, n5171, n5172,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5183, n5184,
         n5185, n5187, n5188, n5190, n5191, n5193, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5214, n5215, n5216, n5217, n5218, n5219, n5222, n5223, n5225,
         n5226, n5227, n5228, n5229, n5230, n5232, n5233, n5234, n5236, n5238,
         n5239, n5240, n5241, n5243, n5244, n5245, n5246, n5247, n5248, n5250,
         n5251, n5253, n5255, n5256, n5257, n5258, n5260, n5261, n5262, n5263,
         n5264, n5267, n5269, n5270, n5271, n5272, n5273, n5275, n5277, n5279,
         n5280, n5282, n5283, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5294, n5295, n5296, n5297, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5307, n5308, n5309, n5310, n5311, n5313, n5316, n5317,
         n5318, n5319, n5321, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5342, n5343, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5365, n5366, n5367, n5368, n5369, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5381, n5382, n5383, n5384, n5385, n5386,
         n5387, n5388, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5407, n5408, n5409, n5411,
         n5412, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5428, n5429, n5430, n5432, n5436, n5437, n5438, n5439,
         n5443, n5444, n5445, n5446, n5448, n5450, n5451, n5452, n5453, n5454,
         n5455, n5457, n5460, n5461, n5462, n5463, n5464, n5467, n5468, n5469,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5483, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5519, n5521, n5522, n5524, n5525, n5526, n5528, n5529,
         n5530, n5532, n5533, n5534, n5536, n5537, n5538, n5539, n5541, n5543,
         n5545, n5546, n5547, n5549, n5551, n5552, n5553, n5554, n5555, n5556,
         n5557, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5568,
         n5569, n5571, n5572, n5574, n5576, n5577, n5578, n5580, n5583, n5584,
         n5586, n5587, n5588, n5589, n5590, n5592, n5593, n5594, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5605, n5606, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5618, n5619, n5620,
         n5622, n5623, n5624, n5627, n5628, n5629, n5630, n5632, n5635, n5637,
         n5638, n5639, n5640, n5641, n5643, n5645, n5646, n5649, n5650, n5651,
         n5653, n5654, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5666, n5667, n5668, n5670, n5671, n5672, n5673, n5674, n5675,
         n5677, n5678, n5679, n5680, n5681, n5682, n5685, n5686, n5688, n5692,
         n5694, n5695, n5696, n5698, n5699, n5700, n5701, n5702, n5703, n5706,
         n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5731, n5733,
         n5735, n5736, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5750,
         n5751, n5752, n5754, n5755, n5757, n5758, n5759, n5760, n5761, n5764,
         n5765, n5766, n5767, n5769, n5770, n5772, n5773, n5774, n5777, n5780,
         n5781, n5783, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5795, n5796, n5799, n5800, n5801, n5803, n5804, n5805, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5819,
         n5820, n5821, n5822, n5823, n5824, n5827, n5828, n5829, n5830, n5831,
         n5832, n5836, n5838, n5840, n5841, n5842, n5843, n5844, n5845, n5847,
         n5848, n5850, n5852, n5853, n5854, n5856, n5857, n5859, n5860, n5861,
         n5863, n5865, n5866, n5867, n5868, n5869, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5895,
         n5896, n5897, n5899, n5900, n5901, n5903, n5905, n5907, n5908, n5909,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5921,
         n5922, n5923, n5924, n5925, n5926, n5928, n5929, n5930, n5932, n5934,
         n5935, n5936, n5938, n5940, n5941, n5942, n5943, n5945, n5946, n5947,
         n5948, n5950, n5951, n5953, n5954, n5955, n5956, n5960, n5961, n5962,
         n5963, n5965, n5966, n5967, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5981, n5983, n5984, n5985, n5986, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5998, n5999, n6000,
         n6001, n6002, n6003, n6005, n6006, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6019, n6020, n6021, n6022, n6023,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6034, n6035, n6036,
         n6037, n6040, n6041, n6042, n6043, n6044, n6046, n6047, n6048, n6049,
         n6050, n6052, n6053, n6054, n6055, n6057, n6058, n6059, n6060, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6071, n6073, n6075,
         n6076, n6077, n6078, n6080, n6081, n6082, n6085, n6086, n6087, n6088,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6099, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6114, n6116, n6118, n6120, n6121, n6122, n6124, n6125, n6126, n6127,
         n6128, n6129, n6130, n6131, n6132, n6134, n6135, n6136, n6137, n6141,
         n6142, n6143, n6144, n6145, n6148, n6149, n6150, n6151, n6153, n6154,
         n6156, n6158, n6159, n6161, n6163, n6164, n6165, n6167, n6168, n6169,
         n6171, n6172, n6175, n6177, n6178, n6180, n6181, n6182, n6183, n6184,
         n6186, n6187, n6188, n6190, n6191, n6192, n6193, n6194, n6195, n6196,
         n6197, n6198, n6201, n6202, n6203, n6204, n6205, n6206, n6208, n6210,
         n6211, n6213, n6214, n6215, n6216, n6217, n6219, n6220, n6221, n6222,
         n6223, n6224, n6226, n6227, n6228, n6230, n6231, n6232, n6233, n6234,
         n6236, n6237, n6238, n6239, n6241, n6243, n6244, n6245, n6247, n6248,
         n6249, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6260,
         n6261, n6262, n6263, n6265, n6266, n6269, n6271, n6272, n6274, n6275,
         n6277, n6278, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6288,
         n6289, n6290, n6292, n6294, n6295, n6296, n6298, n6299, n6300, n6301,
         n6302, n6304, n6306, n6307, n6308, n6309, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6325,
         n6326, n6327, n6329, n6331, n6332, n6333, n6334, n6335, n6336, n6337,
         n6338, n6339, n6340, n6341, n6342, n6343, n6346, n6347, n6349, n6350,
         n6351, n6352, n6353, n6354, n6357, n6359, n6361, n6362, n6363, n6364,
         n6365, n6367, n6369, n6370, n6372, n6373, n6374, n6375, n6376, n6377,
         n6378, n6379, n6380, n6381, n6382, n6384, n6385, n6386, n6387, n6391,
         n6392, n6393, n6394, n6396, n6398, n6399, n6401, n6402, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6412, n6414, n6415, n6416, n6417,
         n6418, n6419, n6420, n6421, n6422, n6424, n6426, n6427, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6438, n6439, n6440, n6441,
         n6442, n6444, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6467, n6468, n6470, n6471, n6472, n6473, n6474, n6476, n6477,
         n6478, n6479, n6480, n6482, n6483, n6485, n6486, n6487, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6497, n6498, n6499, n6500, n6501,
         n6503, n6504, n6505, n6506, n6509, n6510, n6511, n6513, n6514, n6515,
         n6516, n6517, n6518, n6520, n6521, n6522, n6524, n6526, n6527, n6528,
         n6530, n6532, n6534, n6535, n6536, n6537, n6539, n6541, n6542, n6545,
         n6546, n6549, n6551, n6554, n6557, n6559, n6561, n6563, n6564, n6568,
         n6569, n6570, n6573, n6574, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6587, n6588, n6591, n6592, n6593, n6594, n6595,
         n6597, n6602, n6603, n6604, n6605, n6607, n6608, n6609, n6610, n6611,
         n6612, n6614, n6615, n6616, n6617, n6619, n6620, n6622, n6623, n6624,
         n6625, n6626, n6627, n6629, n6631, n6632, n6633, n6634, n6635, n6636,
         n6637, n6640, n6642, n6643, n6644, n6645, n6647, n6648, n6649, n6650,
         n6651, n6652, n6656, n6657, n6660, n6661, n6662, n6663, n6665, n6666,
         n6667, n6668, n6669, n6671, n6672, n6673, n6674, n6678, n6679, n6680,
         n6681, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6694, n6695, n6696, n6697, n6700, n6702, n6703, n6704, n6705, n6706,
         n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717,
         n6718, n6719, n6720, n6721, n6722, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6733, n6734, n6735, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6748, n6749, n6750, n6751, n6754, n6755,
         n6756, n6757, n6758, n6760, n6761, n6762, n6763, n6764, n6765, n6766,
         n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6807, n6808, n6809, n6810, n6811, n6812,
         n6814, n6815, n6816, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6839, n6841, n6843, n6844, n6845, n6846, n6847, n6848, n6850, n6851,
         n6852, n6853, n6854, n6856, n6857, n6858, n6859, n6860, n6862, n6863,
         n6864, n6865, n6867, n6868, n6869, n6870, n6872, n6873, n6874, n6876,
         n6877, n6878, n6879, n6880, n6881, n6883, n6885, n6886, n6887, n6888,
         n6889, n6891, n6893, n6895, n6896, n6898, n6899, n6900, n6902, n6903,
         n6904, n6905, n6906, n6907, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6920, n6921, n6924, n6925, n6926, n6927,
         n6928, n6929, n6930, n6932, n6933, n6935, n6936, n6937, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6947, n6949, n6950, n6951, n6952,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6976, n6977, n6978, n6980, n6981, n6983, n6984, n6985, n6986, n6987,
         n6988, n6989, n6991, n6992, n6994, n6995, n6996, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7018, n7020, n7021, n7024, n7025, n7026, n7027,
         n7028, n7029, n7030, n7031, n7032, n7033, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7043, n7044, n7046, n7048, n7049, n7051, n7052,
         n7053, n7054, n7055, n7056, n7058, n7059, n7060, n7061, n7063, n7064,
         n7065, n7068, n7070, n7071, n7073, n7074, n7077, n7078, n7080, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7094, n7095, n7096, n7098, n7099, n7100, n7101, n7102, n7103, n7106,
         n7107, n7108, n7110, n7111, n7112, n7113, n7114, n7116, n7118, n7119,
         n7120, n7122, n7123, n7124, n7125, n7126, n7128, n7129, n7130, n7131,
         n7132, n7134, n7135, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7151, n7154, n7156, n7157,
         n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7167, n7168,
         n7169, n7170, n7171, n7172, n7174, n7175, n7177, n7178, n7179, n7180,
         n7181, n7185, n7186, n7187, n7189, n7190, n7191, n7192, n7193, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7206,
         n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217,
         n7218, n7219, n7220, n7221, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7233, n7234, n7235, n7236, n7238, n7239, n7241,
         n7246, n7247, n7248, n7249, n7250, n7252, n7253, n7254, n7256, n7257,
         n7258, n7259, n7262, n7263, n7264, n7266, n7267, n7268, n7269, n7270,
         n7272, n7273, n7274, n7275, n7276, n7277, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7289, n7290, n7291, n7292, n7294,
         n7295, n7296, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7308, n7309, n7310, n7311, n7313, n7314, n7315, n7316, n7317,
         n7319, n7320, n7321, n7323, n7324, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7343, n7344, n7345, n7346, n7347, n7349, n7350, n7351, n7352,
         n7353, n7354, n7356, n7357, n7358, n7359, n7360, n7362, n7364, n7366,
         n7367, n7368, n7369, n7370, n7373, n7374, n7375, n7376, n7378, n7381,
         n7382, n7383, n7384, n7385, n7386, n7388, n7389, n7391, n7392, n7393,
         n7394, n7395, n7396, n7400, n7401, n7404, n7406, n7407, n7409, n7410,
         n7411, n7413, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7426, n7427, n7428, n7429, n7430, n7431, n7433, n7434, n7435, n7436,
         n7437, n7439, n7440, n7442, n7443, n7444, n7446, n7447, n7450, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7466, n7468, n7469, n7471, n7472, n7473, n7474, n7475,
         n7477, n7478, n7479, n7480, n7481, n7483, n7484, n7485, n7486, n7487,
         n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7498,
         n7499, n7500, n7501, n7502, n7504, n7505, n7506, n7507, n7508, n7509,
         n7511, n7512, n7513, n7515, n7516, n7517, n7518, n7521, n7522, n7523,
         n7526, n7527, n7528, n7529, n7530, n7532, n7533, n7534, n7535, n7536,
         n7537, n7539, n7540, n7541, n7543, n7544, n7545, n7546, n7547, n7548,
         n7550, n7551, n7554, n7555, n7556, n7557, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7568, n7569, n7570, n7571, n7572, n7573,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7587, n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596,
         n7597, n7598, n7599, n7600, n7601, n7602, n7605, n7607, n7608, n7609,
         n7610, n7613, n7614, n7616, n7617, n7618, n7619, n7620, n7622, n7623,
         n7624, n7626, n7627, n7628, n7629, n7630, n7631, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7642, n7643, n7644, n7645, n7646,
         n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7657,
         n7658, n7659, n7660, n7661, n7662, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7674, n7675, n7676, n7677, n7680, n7682, n7683,
         n7685, n7686, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7699, n7700, n7702, n7704, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7720,
         n7721, n7722, n7724, n7725, n7726, n7728, n7729, n7730, n7732, n7733,
         n7735, n7736, n7737, n7739, n7740, n7741, n7742, n7743, n7746, n7747,
         n7748, n7749, n7750, n7751, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7768, n7769, n7770,
         n7772, n7773, n7774, n7775, n7776, n7777, n7780, n7782, n7783, n7784,
         n7785, n7786, n7788, n7789, n7790, n7791, n7792, n7793, n7795, n7796,
         n7797, n7798, n7799, n7800, n7802, n7803, n7804, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7820, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7860, n7861, n7862, n7864, n7865, n7866,
         n7867, n7868, n7870, n7871, n7872, n7873, n7875, n7876, n7877, n7878,
         n7881, n7882, n7883, n7884, n7886, n7888, n7889, n7890, n7892, n7893,
         n7894, n7895, n7896, n7898, n7899, n7900, n7902, n7903, n7904, n7905,
         n7906, n7907, n7909, n7911, n7912, n7913, n7914, n7915, n7916, n7918,
         n7919, n7920, n7922, n7923, n7924, n7925, n7926, n7927, n7929, n7930,
         n7931, n7932, n7933, n7935, n7936, n7938, n7939, n7943, n7944, n7945,
         n7946, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956,
         n7957, n7958, n7959, n7960, n7962, n7963, n7964, n7965, n7966, n7967,
         n7968, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7978, n7979,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8018, n8019, n8020, n8021, n8023, n8024, n8026, n8027,
         n8029, n8030, n8031, n8033, n8034, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8045, n8047, n8050, n8052, n8053, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8072, n8074, n8075, n8076, n8077, n8078,
         n8080, n8081, n8082, n8084, n8086, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8100, n8102, n8103, n8104, n8105, n8106, n8107,
         n8109, n8110, n8111, n8112, n8113, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8123, n8125, n8126, n8127, n8128, n8129, n8130, n8131,
         n8132, n8133, n8134, n8135, n8137, n8139, n8141, n8142, n8144, n8145,
         n8146, n8147, n8148, n8151, n8152, n8153, n8154, n8157, n8158, n8159,
         n8160, n8161, n8162, n8164, n8165, n8167, n8168, n8169, n8170, n8171,
         n8172, n8173, n8174, n8176, n8177, n8178, n8179, n8180, n8183, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8193, n8194, n8195, n8196,
         n8197, n8198, n8201, n8203, n8204, n8206, n8207, n8208, n8209, n8211,
         n8212, n8214, n8215, n8216, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8233, n8234, n8235, n8237,
         n8238, n8240, n8241, n8243, n8244, n8245, n8246, n8248, n8249, n8250,
         n8251, n8252, n8254, n8257, n8258, n8259, n8261, n8263, n8264, n8266,
         n8267, n8268, n8269, n8271, n8272, n8274, n8275, n8277, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8287, n8289, n8290, n8292, n8294,
         n8295, n8296, n8297, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8310, n8311, n8312, n8313, n8315, n8316, n8317,
         n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327,
         n8328, n8329, n8331, n8332, n8333, n8334, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8346, n8347, n8348, n8350, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8361, n8362, n8363, n8364,
         n8365, n8367, n8368, n8369, n8370, n8371, n8373, n8375, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8385, n8386, n8388, n8389, n8390,
         n8391, n8393, n8394, n8396, n8397, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8420, n8421, n8422, n8423, n8424, n8426,
         n8427, n8428, n8429, n8430, n8431, n8433, n8434, n8435, n8436, n8437,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8449,
         n8450, n8452, n8453, n8454, n8455, n8456, n8458, n8459, n8460, n8461,
         n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8471, n8472,
         n8473, n8474, n8475, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8491, n8492, n8494, n8497,
         n8498, n8499, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8512, n8513, n8515, n8517, n8518, n8520, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8531, n8532, n8533, n8534,
         n8535, n8536, n8539, n8541, n8542, n8543, n8544, n8545, n8546, n8547,
         n8549, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8560, n8561,
         n8563, n8564, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8574,
         n8575, n8576, n8577, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8597,
         n8598, n8599, n8601, n8602, n8604, n8605, n8606, n8608, n8609, n8610,
         n8611, n8613, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8658,
         n8659, n8660, n8661, n8662, n8664, n8665, n8666, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8688, n8689, n8690, n8691,
         n8692, n8693, n8694, n8695, n8696, n8698, n8699, n8700, n8701, n8703,
         n8704, n8707, n8709, n8710, n8711, n8712, n8714, n8716, n8717, n8718,
         n8719, n8720, n8722, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741,
         n8742, n8743, n8744, n8745, n8746, n8750, n8751, n8752, n8753, n8755,
         n8756, n8758, n8759, n8760, n8761, n8763, n8764, n8765, n8766, n8767,
         n8768, n8769, n8770, n8772, n8773, n8774, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8785, n8787, n8788, n8789, n8790, n8792,
         n8793, n8794, n8796, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8815, n8817,
         n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827,
         n8828, n8829, n8830, n8831, n8832, n8834, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8854, n8855, n8856, n8857, n8858, n8859, n8862,
         n8863, n8864, n8865, n8866, n8867, n8869, n8870, n8873, n8874, n8875,
         n8876, n8878, n8879, n8881, n8882, n8884, n8887, n8888, n8890, n8892,
         n8893, n8894, n8895, n8897, n8899, n8900, n8901, n8903, n8904, n8906,
         n8907, n8908, n8909, n8910, n8914, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8926, n8927, n8928, n8930, n8931, n8933, n8935, n8936,
         n8937, n8938, n8940, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8962, n8963, n8964, n8965, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8976, n8977, n8978, n8979, n8980, n8983, n8984, n8985,
         n8986, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8998, n8999, n9000, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9027, n9028, n9029, n9031, n9032,
         n9033, n9035, n9036, n9037, n9038, n9040, n9042, n9044, n9046, n9048,
         n9049, n9050, n9052, n9053, n9054, n9057, n9060, n9062, n9063, n9065,
         n9066, n9067, n9069, n9070, n9071, n9072, n9073, n9075, n9076, n9077,
         n9078, n9079, n9081, n9082, n9083, n9085, n9086, n9087, n9088, n9090,
         n9092, n9093, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9107, n9108, n9110, n9111, n9112, n9113, n9114, n9115,
         n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9136, n9137, n9138, n9139, n9140,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9156, n9158, n9159, n9160, n9161, n9163, n9166, n9167,
         n9168, n9169, n9170, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9180, n9181, n9183, n9184, n9185, n9186, n9187, n9189, n9190, n9191,
         n9193, n9194, n9195, n9196, n9197, n9199, n9201, n9202, n9203, n9206,
         n9207, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217,
         n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227,
         n9229, n9230, n9231, n9232, n9233, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9259, n9260,
         n9261, n9263, n9264, n9266, n9267, n9268, n9269, n9271, n9272, n9273,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9285,
         n9286, n9287, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317,
         n9318, n9319, n9320, n9321, n9323, n9325, n9326, n9328, n9329, n9331,
         n9332, n9333, n9334, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9346, n9347, n9348, n9349, n9350, n9352, n9354, n9355, n9356,
         n9357, n9358, n9359, n9361, n9362, n9363, n9364, n9365, n9366, n9367,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9404, n9405, n9406, n9407, n9408, n9410, n9412,
         n9415, n9416, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427,
         n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437,
         n9438, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9449,
         n9451, n9453, n9454, n9455, n9456, n9457, n9459, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9481, n9482, n9483, n9484,
         n9485, n9487, n9490, n9491, n9492, n9493, n9494, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9506, n9508, n9509, n9510,
         n9511, n9512, n9514, n9515, n9516, n9517, n9518, n9521, n9522, n9523,
         n9524, n9525, n9526, n9528, n9529, n9530, n9531, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9551, n9552, n9554, n9555, n9557, n9558, n9559,
         n9560, n9562, n9563, n9564, n9565, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9576, n9577, n9578, n9579, n9580, n9581, n9583, n9584,
         n9585, n9586, n9590, n9591, n9592, n9594, n9597, n9598, n9599, n9601,
         n9602, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9632, n9634, n9636, n9637, n9638,
         n9640, n9641, n9642, n9643, n9645, n9647, n9649, n9651, n9652, n9653,
         n9654, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9670, n9671, n9672, n9675, n9677, n9678, n9679,
         n9680, n9681, n9684, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9694, n9695, n9696, n9697, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9710, n9711, n9712, n9713, n9714, n9715,
         n9717, n9718, n9719, n9720, n9721, n9722, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9740,
         n9741, n9742, n9743, n9744, n9745, n9747, n9748, n9749, n9751, n9752,
         n9753, n9754, n9755, n9757, n9758, n9759, n9761, n9762, n9763, n9764,
         n9765, n9767, n9768, n9769, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9781, n9782, n9783, n9784, n9785, n9786, n9788,
         n9789, n9790, n9791, n9792, n9793, n9795, n9796, n9797, n9798, n9799,
         n9801, n9803, n9805, n9807, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9822, n9823, n9824, n9825, n9826,
         n9827, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837,
         n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847,
         n9848, n9849, n9850, n9851, n9853, n9855, n9856, n9857, n9858, n9859,
         n9860, n9862, n9863, n9864, n9865, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9900, n9901, n9902, n9903, n9904,
         n9906, n9907, n9908, n9909, n9910, n9911, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9959, n9960,
         n9961, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9971, n9972,
         n9974, n9975, n9977, n9978, n9980, n9981, n9982, n9983, n9984, n9986,
         n9987, n9988, n9989, n9990, n9991, n9993, n9994, n9995, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10038, n10039, n10040, n10041, n10042,
         n10044, n10045, n10046, n10047, n10049, n10050, n10051, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10069, n10071,
         n10072, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10085, n10086, n10087, n10088, n10090,
         n10091, n10093, n10094, n10096, n10097, n10098, n10099, n10100,
         n10102, n10103, n10104, n10106, n10107, n10108, n10109, n10111,
         n10112, n10113, n10114, n10115, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10131, n10132, n10133, n10134, n10135, n10137, n10138,
         n10140, n10141, n10142, n10143, n10144, n10146, n10147, n10148,
         n10149, n10151, n10152, n10153, n10155, n10156, n10157, n10158,
         n10159, n10160, n10161, n10162, n10163, n10164, n10166, n10167,
         n10169, n10171, n10172, n10173, n10174, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10207, n10208, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10219, n10220, n10221, n10222,
         n10223, n10224, n10225, n10226, n10228, n10229, n10230, n10232,
         n10234, n10235, n10237, n10238, n10239, n10240, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10255,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10288, n10289,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10300,
         n10301, n10303, n10304, n10306, n10307, n10309, n10310, n10311,
         n10312, n10314, n10315, n10316, n10317, n10319, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10331,
         n10332, n10333, n10334, n10335, n10337, n10338, n10339, n10341,
         n10342, n10343, n10344, n10346, n10347, n10348, n10349, n10350,
         n10351, n10352, n10353, n10354, n10356, n10357, n10359, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10373, n10375, n10378, n10379, n10382, n10384,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10400, n10402, n10403,
         n10404, n10405, n10407, n10408, n10411, n10412, n10413, n10414,
         n10415, n10416, n10417, n10418, n10419, n10420, n10421, n10422,
         n10423, n10425, n10426, n10427, n10428, n10429, n10430, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10455, n10456, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10484, n10485, n10486,
         n10487, n10488, n10489, n10490, n10491, n10492, n10493, n10496,
         n10497, n10498, n10499, n10500, n10501, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10514,
         n10515, n10516, n10519, n10520, n10521, n10522, n10523, n10524,
         n10525, n10526, n10527, n10528, n10530, n10532, n10533, n10534,
         n10535, n10536, n10537, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10571, n10572, n10574, n10575, n10576, n10577, n10579, n10580,
         n10581, n10582, n10583, n10585, n10586, n10587, n10588, n10590,
         n10591, n10592, n10593, n10594, n10595, n10596, n10597, n10598,
         n10599, n10600, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10613, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10627, n10628,
         n10629, n10630, n10631, n10632, n10633, n10634, n10635, n10636,
         n10638, n10640, n10641, n10642, n10643, n10644, n10645, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10657,
         n10658, n10659, n10661, n10662, n10663, n10664, n10665, n10667,
         n10668, n10669, n10671, n10673, n10674, n10676, n10677, n10678,
         n10679, n10680, n10682, n10683, n10684, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10694, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10706, n10707,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10730, n10731, n10732, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10742, n10744, n10745,
         n10746, n10747, n10748, n10750, n10751, n10752, n10753, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10770, n10771, n10772,
         n10773, n10774, n10775, n10776, n10778, n10779, n10780, n10781,
         n10782, n10783, n10785, n10786, n10788, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10827, n10828,
         n10829, n10830, n10831, n10832, n10833, n10834, n10835, n10836,
         n10837, n10838, n10839, n10840, n10841, n10843, n10844, n10845,
         n10847, n10848, n10849, n10850, n10851, n10852, n10853, n10855,
         n10856, n10859, n10860, n10861, n10862, n10863, n10864, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10879, n10880, n10881, n10882, n10883,
         n10884, n10886, n10887, n10888, n10889, n10890, n10892, n10893,
         n10895, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10944, n10945, n10946,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10960, n10961, n10962, n10963, n10965, n10966,
         n10967, n10969, n10970, n10972, n10973, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10986,
         n10987, n10988, n10989, n10990, n10991, n10993, n10994, n10995,
         n10997, n10998, n10999, n11001, n11002, n11003, n11004, n11005,
         n11007, n11008, n11009, n11010, n11011, n11012, n11013, n11014,
         n11015, n11016, n11017, n11018, n11020, n11021, n11022, n11023,
         n11025, n11026, n11027, n11028, n11029, n11030, n11032, n11033,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11070,
         n11071, n11072, n11073, n11074, n11075, n11076, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11095, n11096, n11097, n11099,
         n11100, n11101, n11103, n11104, n11105, n11106, n11108, n11109,
         n11110, n11111, n11113, n11114, n11115, n11116, n11117, n11118,
         n11119, n11120, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11142, n11143, n11144,
         n11145, n11146, n11147, n11150, n11151, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11162, n11163, n11164,
         n11167, n11168, n11170, n11171, n11172, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11200, n11201, n11203, n11204, n11205, n11206,
         n11207, n11208, n11211, n11212, n11213, n11215, n11217, n11218,
         n11219, n11220, n11221, n11223, n11224, n11225, n11226, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11311, n11314, n11315, n11316, n11319, n11320, n11321, n11323,
         n11324, n11325, n11326, n11327, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11340, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11352,
         n11353, n11354, n11355, n11356, n11357, n11359, n11360, n11361,
         n11362, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11375, n11376, n11377, n11378, n11380,
         n11382, n11383, n11384, n11385, n11386, n11388, n11389, n11390,
         n11391, n11392, n11393, n11394, n11395, n11396, n11398, n11400,
         n11401, n11402, n11403, n11404, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11444, n11445,
         n11447, n11448, n11450, n11451, n11452, n11453, n11454, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11507, n11508, n11509,
         n11511, n11513, n11514, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11527, n11529, n11530,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11546, n11548, n11549, n11550,
         n11551, n11552, n11553, n11554, n11556, n11557, n11558, n11559,
         n11560, n11561, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11595,
         n11596, n11599, n11600, n11601, n11602, n11604, n11605, n11606,
         n11608, n11609, n11610, n11611, n11613, n11615, n11616, n11617,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11632, n11633, n11635, n11636,
         n11637, n11638, n11639, n11640, n11642, n11643, n11644, n11645,
         n11646, n11648, n11649, n11650, n11652, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11684, n11685, n11686, n11687, n11688, n11689, n11691,
         n11692, n11693, n11695, n11696, n11697, n11700, n11701, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11741, n11742, n11743, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11765,
         n11766, n11767, n11768, n11770, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11781, n11782, n11783, n11784, n11785,
         n11786, n11788, n11790, n11791, n11792, n11794, n11795, n11796,
         n11797, n11798, n11800, n11801, n11802, n11803, n11804, n11806,
         n11807, n11808, n11809, n11810, n11811, n11812, n11814, n11815,
         n11816, n11818, n11819, n11820, n11821, n11822, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11893,
         n11894, n11895, n11896, n11898, n11899, n11900, n11901, n11903,
         n11904, n11908, n11909, n11910, n11912, n11913, n11914, n11915,
         n11916, n11918, n11919, n11921, n11923, n11924, n11925, n11927,
         n11928, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11939, n11940, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11951, n11952, n11953, n11954, n11955, n11956,
         n11959, n11960, n11961, n11962, n11963, n11964, n11965, n11966,
         n11967, n11968, n11970, n11971, n11972, n11973, n11976, n11977,
         n11978, n11980, n11981, n11983, n11984, n11985, n11986, n11989,
         n11990, n11991, n11992, n11993, n11994, n11997, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12015, n12016, n12017,
         n12018, n12020, n12021, n12022, n12023, n12024, n12026, n12027,
         n12028, n12030, n12031, n12032, n12033, n12035, n12036, n12038,
         n12040, n12041, n12042, n12043, n12044, n12045, n12047, n12048,
         n12052, n12054, n12055, n12059, n12060, n12061, n12063, n12064,
         n12065, n12068, n12069, n12071, n12072, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12176, n12177, n12178, n12179, n12180, n12181, n12182,
         n12183, n12184, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, N28617, N28616, N28615, N28613, N28612, N28611, N28610,
         N28609, N28608, N28607, N28606, N28598, N28597, N28590, N28589,
         N28588, N28582, N28581, N28580, N28579, N28576, N28575, N28574,
         N28573, N28572, N28571, N28570, N28562, N28561, N28553, N28552,
         N28545, N28544, N28543, N28536, N28535, N28534, N28527, N28526,
         N28525, N28519, N28518, N28517, N28516, N28511, N28510, N28509,
         N28508, N28507, N28504, N28503, N28502, N28501, N28500, N28499,
         N28498, N28490, N28489, N28481, N28480, N28472, N28471, N28463,
         N28462, N28454, N28453, N28446, N28445, N28444, N28437, N28436,
         N28435, N28428, N28427, N28426, N28419, N28418, N28417, N28410,
         N28409, N28408, N28401, N28400, N28399, N28393, N28392, N28391,
         N28390, N28384, N28383, N28382, N28381, N28376, N28375, N28374,
         N28373, N28372, N28367, N28366, N28365, N28364, N28363, N28360,
         N28359, N28358, N28357, N28356, N28355, N28354, N28346, N28345,
         N28337, N28336, N28328, N28327, N28319, N28318, N28310, N28309,
         N28301, N28300, N28292, N28291, N28283, N28282, N28274, N28273,
         N28265, N28264, N28256, N28255, N28248, N28247, N28246, N28239,
         N28238, N28237, N28230, N28229, N28228, N28221, N28220, N28219,
         N28212, N28211, N28210, N28203, N28202, N28201, N28194, N28193,
         N28192, N28185, N28184, N28183, N28176, N28175, N28174, N28167,
         N28166, N28165, N28158, N28157, N28156, N28150, N28149, N28148,
         N28147, N28141, N28140, N28139, N28138, N28132, N28131, N28130,
         N28129, N28123, N28122, N28121, N28120, N28114, N28113, N28112,
         N28111, N28106, N28105, N28104, N28103, N28102, N28097, N28096,
         N28095, N28094, N28093, N28088, N28087, N28086, N28085, N28084,
         N28080, N28079, N28078, N28077, N28076, N28075, N28071, N28070,
         N28069, N28068, N28067, N28066, N28058, N28057, N28049, N28048,
         N28040, N28039, N28031, N28030, N28022, N28021, N28013, N28012,
         N28004, N28003, N27995, N27994, N27986, N27985, N27977, N27976,
         N27968, N27967, N27959, N27958, N27950, N27949, N27941, N27940,
         N27932, N27931, N27923, N27922, N27914, N27913, N27905, N27904,
         N27896, N27895, N27887, N27886, N27878, N27877, N27869, N27868,
         N27860, N27859, N27851, N27850, N27843, N27842, N27841, N27834,
         N27833, N27832, N27825, N27824, N27823, N27816, N27815, N27814,
         N27807, N27806, N27805, N27798, N27797, N27796, N27789, N27788,
         N27787, N27780, N27779, N27778, N27771, N27770, N27769, N27762,
         N27761, N27760, N27753, N27752, N27751, N27744, N27743, N27742,
         N27735, N27734, N27733, N27726, N27725, N27724, N27717, N27716,
         N27715, N27708, N27707, N27706, N27699, N27698, N27697, N27690,
         N27689, N27688, N27681, N27680, N27679, N27672, N27671, N27670,
         N27664, N27663, N27662, N27661, N27655, N27654, N27653, N27652,
         N27646, N27645, N27644, N27643, N27637, N27636, N27635, N27634,
         N27628, N27627, N27626, N27625, N27619, N27618, N27617, N27616,
         N27610, N27609, N27608, N27607, N27601, N27600, N27599, N27598,
         N27592, N27591, N27590, N27589, N27583, N27582, N27581, N27580,
         N27574, N27573, N27572, N27571, N27565, N27564, N27563, N27562,
         N27557, N27556, N27555, N27554, N27553, N27548, N27547, N27546,
         N27545, N27544, N27539, N27538, N27537, N27536, N27535, N27530,
         N27529, N27528, N27527, N27526, N27521, N27520, N27519, N27518,
         N27517, N27513, N27512, N27511, N27510, N27509, N27508, N27504,
         N27503, N27502, N27501, N27500, N27499, N27495, N27494, N27493,
         N27492, N27491, N27490, N27482, N27481, N27473, N27472, N27464,
         N27463, N27455, N27454, N27446, N27445, N27437, N27436, N27428,
         N27427, N27419, N27418, N27410, N27409, N27401, N27400, N27392,
         N27391, N27383, N27382, N27374, N27373, N27365, N27364, N27356,
         N27355, N27347, N27346, N27338, N27337, N27329, N27328, N27320,
         N27319, N27311, N27310, N27302, N27301, N27293, N27292, N27284,
         N27283, N27275, N27274, N27266, N27265, N27257, N27256, N27248,
         N27247, N27239, N27238, N27230, N27229, N27221, N27220, N27212,
         N27211, N27203, N27202, N27194, N27193, N27185, N27184, N27176,
         N27175, N27167, N27166, N27158, N27157, N27149, N27148, N27140,
         N27139, N27131, N27130, N27122, N27121, N27113, N27112, N29417,
         N29416, N29415, N29414, N3855, N29401, N29400, N29399, N4664, N29405,
         N29404, N29403, \lt_82/A[5] , \lt_82/A[4] , \sub_183/carry[8] ,
         \sub_183/carry[7] , \sub_183/carry[6] , \sub_183/carry[5] ,
         \sub_183/carry[4] , \sub_183/carry[3] ,
         \add_1_root_add_115_2/carry[11] , \add_1_root_add_115_2/carry[10] ,
         \add_114/carry[11] , \add_114/carry[10] ,
         \add_1_root_add_89_2/carry[11] , \add_1_root_add_89_2/carry[10] ,
         \add_0_root_add_0_root_add_129_2/carry[11] ,
         \add_0_root_add_0_root_add_129_2/carry[10] ,
         \add_0_root_add_0_root_add_129_2/carry[9] ,
         \add_0_root_add_0_root_add_129_2/carry[8] ,
         \add_0_root_add_0_root_add_129_2/carry[7] ,
         \add_0_root_add_0_root_add_129_2/carry[6] ,
         \add_0_root_add_0_root_add_129_2/carry[5] ,
         \add_0_root_add_0_root_add_129_2/carry[4] ,
         \add_0_root_add_1_root_add_130_3/carry[11] ,
         \add_0_root_add_1_root_add_130_3/carry[10] ,
         \add_0_root_add_1_root_add_130_3/carry[9] ,
         \add_0_root_add_1_root_add_130_3/carry[8] ,
         \add_0_root_add_1_root_add_130_3/carry[7] ,
         \add_0_root_add_1_root_add_130_3/carry[6] ,
         \add_0_root_add_1_root_add_130_3/carry[5] ,
         \add_0_root_add_1_root_add_130_3/carry[4] ,
         \add_1_root_add_158_3/carry[11] , \add_1_root_add_158_3/carry[10] ,
         \add_157_2/carry[11] , \add_157_2/carry[10] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[5] ,
         \add_1_root_add_86_root_add_255_countones_143/carry[6] ,
         \add_2_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_2_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_2_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_2_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_2_root_add_86_root_add_255_countones_143/carry[5] ,
         \add_3_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_3_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_3_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_3_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_3_root_add_86_root_add_255_countones_143/carry[5] ,
         \add_4_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_4_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_4_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_4_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_4_root_add_86_root_add_255_countones_143/carry[5] ,
         \add_11_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_11_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_11_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_8_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_8_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_8_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_8_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_18_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_18_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_18_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_27_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_27_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_58_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_19_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_19_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_19_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_5_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_5_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_5_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_5_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_12_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_12_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_12_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_26_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_26_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_54_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_49_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_47_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_38_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_38_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_65_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_73_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_37_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_37_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_66_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_76_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_28_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_28_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_46_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_55_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_25_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_25_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_63_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_52_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_24_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_24_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_56_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_51_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_21_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_21_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_67_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_60_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_17_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_17_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_17_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_32_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_32_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_79_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_72_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_36_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_36_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_80_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_75_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_9_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_9_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_9_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_9_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_10_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_10_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_10_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_35_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_35_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_68_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_71_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_31_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_31_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_44_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_43_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_20_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_20_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_20_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_41_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_41_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_42_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_53_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_7_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_7_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_7_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_7_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_16_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_16_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_16_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_34_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_34_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_70_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_69_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_33_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_33_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_78_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_62_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_14_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_14_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_14_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_22_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_22_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_57_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_48_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_29_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_29_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_45_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_59_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_6_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_6_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_6_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_6_root_add_86_root_add_255_countones_143/carry[4] ,
         \add_15_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_15_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_15_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_39_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_39_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_64_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_77_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_40_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_40_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_83_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_82_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_13_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_13_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_13_root_add_86_root_add_255_countones_143/carry[3] ,
         \add_23_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_23_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_74_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_50_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_30_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_30_root_add_86_root_add_255_countones_143/carry[2] ,
         \add_81_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_61_root_add_86_root_add_255_countones_143/carry[1] ,
         \add_0_root_add_1_root_add_98_3/carry[11] ,
         \add_0_root_add_1_root_add_98_3/carry[10] ,
         \add_0_root_add_1_root_add_98_3/carry[9] ,
         \add_0_root_add_1_root_add_98_3/carry[8] ,
         \add_0_root_add_1_root_add_98_3/carry[7] ,
         \add_0_root_add_1_root_add_98_3/carry[6] ,
         \add_0_root_add_1_root_add_98_3/carry[5] ,
         \add_0_root_add_1_root_add_98_3/carry[4] ,
         \add_0_root_add_1_root_add_98_3/A[3] ,
         \add_0_root_add_1_root_add_98_3/A[4] ,
         \add_0_root_add_1_root_add_98_3/A[5] ,
         \add_0_root_add_1_root_add_98_3/A[6] ,
         \add_0_root_add_1_root_add_98_3/A[7] ,
         \add_0_root_add_1_root_add_98_3/A[8] ,
         \add_0_root_add_1_root_add_98_3/A[9] ,
         \add_0_root_add_1_root_add_98_3/A[10] ,
         \add_0_root_add_1_root_add_98_3/A[11] ,
         \add_0_root_add_0_root_add_97_2/carry[11] ,
         \add_0_root_add_0_root_add_97_2/carry[10] ,
         \add_0_root_add_0_root_add_97_2/carry[9] ,
         \add_0_root_add_0_root_add_97_2/carry[8] ,
         \add_0_root_add_0_root_add_97_2/carry[7] ,
         \add_0_root_add_0_root_add_97_2/carry[6] ,
         \add_0_root_add_0_root_add_97_2/carry[5] ,
         \add_0_root_add_0_root_add_97_2/carry[4] , \add_88_aco/carry[11] ,
         \add_88_aco/carry[10] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n824,
         n825, n826, n827, n828, n829, n830, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n855, n856, n857, n858, n859, n860,
         n861, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3582, n3586, n3587, n3618, n3619, n3621, n3650,
         n3653, n3659, n3660, n3664, n3665, n3668, n3672, n3675, n3678, n3679,
         n3681, n3684, n3692, n3699, n3700, n3708, n3712, n3715, n3717, n3719,
         n3721, n3723, n3725, n3728, n3730, n3732, n3734, n3736, n3738, n3740,
         n3742, n3744, n3746, n3748, n3751, n3753, n3755, n3757, n3759, n3761,
         n3764, n3766, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3795, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3826, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4195, n4196, n4199, n4201,
         n4203, n4205, n4207, n4209, n4210, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4238, n4239, n4243, n4244, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4255, n4256, n4257,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4326, n4328, n4330, n4331,
         n4334, n4338, n4339, n4342, n4346, n4347, n4352, n4357, n4361, n4365,
         n4366, n4368, n4369, n4373, n4374, n4376, n4383, n4384, n4392, n4393,
         n4396, n4397, n4404, n4405, n4406, n4408, n4411, n4416, n4419, n4421,
         n4423, n4426, n4427, n4436, n4437, n4438, n4439, n4441, n4444, n4450,
         n4451, n4457, n4459, n4462, n4464, n4470, n4471, n4481, n4491, n4493,
         n4497, n4503, n4506, n4510, n4512, n4514, n4523, n4524, n4530, n4549,
         n4551, n4552, n4561, n4568, n4572, n4575, n4576, n4580, n4587, n4590,
         n4595, n4604, n4608, n4619, n4628, n4633, n4635, n4640, n4646, n4649,
         n4653, n4656, n4663, n4668, n4675, n4677, n4681, n4683, n4689, n4691,
         n4692, n4693, n4698, n4703, n4711, n4719, n4725, n4727, n4735, n4742,
         n4745, n4746, n4747, n4751, n4754, n4766, n4767, n4771, n4776, n4789,
         n4793, n4816, n4819, n4827, n4832, n4835, n4844, n4847, n4854, n4858,
         n4866, n4871, n4881, n4886, n4889, n4890, n4894, n4895, n4900, n4901,
         n4902, n4913, n4915, n4922, n4939, n4941, n4944, n4946, n4948, n4949,
         n4951, n4954, n4957, n4958, n4959, n4962, n4965, n4966, n4973, n4974,
         n4976, n4980, n4984, n4998, n4999, n5003, n5034, n5035, n5043, n5044,
         n5046, n5049, n5052, n5060, n5061, n5063, n5068, n5071, n5079, n5093,
         n5096, n5098, n5101, n5104, n5106, n5110, n5113, n5118, n5124, n5126,
         n5129, n5136, n5140, n5142, n5145, n5146, n5152, n5156, n5164, n5165,
         n5168, n5173, n5182, n5186, n5189, n5192, n5194, n5203, n5204, n5205,
         n5213, n5220, n5221, n5224, n5231, n5235, n5237, n5242, n5249, n5252,
         n5254, n5259, n5265, n5266, n5268, n5274, n5276, n5278, n5281, n5284,
         n5293, n5298, n5306, n5312, n5314, n5315, n5320, n5322, n5341, n5344,
         n5354, n5355, n5364, n5370, n5380, n5389, n5397, n5405, n5406, n5410,
         n5413, n5414, n5426, n5427, n5431, n5433, n5434, n5435, n5440, n5441,
         n5442, n5447, n5449, n5456, n5458, n5459, n5465, n5466, n5470, n5482,
         n5484, n5494, n5495, n5506, n5518, n5520, n5523, n5527, n5531, n5535,
         n5540, n5542, n5544, n5548, n5550, n5558, n5567, n5570, n5573, n5575,
         n5579, n5581, n5582, n5585, n5591, n5595, n5604, n5607, n5617, n5621,
         n5625, n5626, n5631, n5633, n5634, n5636, n5642, n5644, n5647, n5648,
         n5652, n5655, n5665, n5669, n5676, n5683, n5684, n5687, n5689, n5690,
         n5691, n5693, n5697, n5704, n5705, n5714, n5715, n5727, n5728, n5729,
         n5730, n5732, n5734, n5737, n5738, n5746, n5747, n5748, n5749, n5753,
         n5756, n5762, n5763, n5768, n5771, n5775, n5776, n5778, n5779, n5782,
         n5784, n5785, n5794, n5797, n5798, n5802, n5806, n5818, n5825, n5826,
         n5833, n5834, n5835, n5837, n5839, n5846, n5849, n5851, n5855, n5858,
         n5862, n5864, n5870, n5894, n5898, n5902, n5904, n5906, n5910, n5920,
         n5927, n5931, n5933, n5937, n5939, n5944, n5949, n5952, n5957, n5958,
         n5959, n5964, n5968, n5979, n5980, n5982, n5987, n5988, n5997, n6004,
         n6007, n6018, n6024, n6025, n6033, n6038, n6039, n6045, n6051, n6056,
         n6061, n6070, n6072, n6074, n6079, n6083, n6084, n6089, n6097, n6098,
         n6100, n6113, n6115, n6117, n6119, n6123, n6133, n6138, n6139, n6140,
         n6146, n6147, n6152, n6155, n6157, n6160, n6162, n6166, n6170, n6173,
         n6174, n6176, n6179, n6185, n6189, n6199, n6200, n6207, n6209, n6212,
         n6218, n6225, n6229, n6235, n6240, n6242, n6246, n6250, n6259, n6264,
         n6267, n6268, n6270, n6273, n6276, n6279, n6287, n6291, n6293, n6297,
         n6303, n6305, n6310, n6324, n6328, n6330, n6344, n6345, n6348, n6355,
         n6356, n6358, n6360, n6366, n6368, n6371, n6383, n6388, n6389, n6390,
         n6395, n6397, n6400, n6403, n6411, n6413, n6423, n6425, n6428, n6437,
         n6443, n6445, n6455, n6466, n6469, n6475, n6481, n6484, n6488, n6496,
         n6502, n6507, n6508, n6512, n6519, n6523, n6525, n6529, n6531, n6533,
         n6538, n6540, n6543, n6544, n6547, n6548, n6550, n6552, n6553, n6555,
         n6556, n6558, n6560, n6562, n6565, n6566, n6567, n6571, n6572, n6575,
         n6576, n6586, n6589, n6590, n6596, n6598, n6599, n6600, n6601, n6606,
         n6613, n6618, n6621, n6628, n6630, n6638, n6639, n6641, n6646, n6653,
         n6654, n6655, n6658, n6659, n6664, n6670, n6675, n6676, n6677, n6682,
         n6683, n6693, n6698, n6699, n6701, n6707, n6723, n6731, n6732, n6736,
         n6737, n6747, n6752, n6753, n6759, n6776, n6777, n6778, n6795, n6805,
         n6806, n6813, n6817, n6818, n6826, n6837, n6838, n6840, n6842, n6849,
         n6855, n6861, n6866, n6871, n6875, n6882, n6884, n6890, n6892, n6894,
         n6897, n6901, n6908, n6919, n6922, n6923, n6931, n6934, n6938, n6946,
         n6948, n6953, n6967, n6975, n6979, n6982, n6990, n6993, n6997, n6998,
         n7006, n7016, n7017, n7019, n7022, n7023, n7034, n7042, n7045, n7047,
         n7050, n7057, n7062, n7066, n7067, n7069, n7072, n7075, n7076, n7079,
         n7081, n7093, n7097, n7104, n7105, n7109, n7115, n7117, n7121, n7127,
         n7133, n7136, n7150, n7152, n7153, n7155, n7166, n7173, n7176, n7182,
         n7183, n7184, n7188, n7194, n7205, n7207, n7222, n7232, n7237, n7240,
         n7242, n7243, n7244, n7245, n7251, n7255, n7260, n7261, n7265, n7271,
         n7278, n7288, n7293, n7297, n7307, n7312, n7318, n7322, n7325, n7342,
         n7348, n7355, n7361, n7363, n7365, n7371, n7372, n7377, n7379, n7380,
         n7387, n7390, n7397, n7398, n7399, n7402, n7403, n7405, n7408, n7412,
         n7414, n7415, n7424, n7425, n7432, n7438, n7441, n7445, n7448, n7449,
         n7451, n7465, n7467, n7470, n7476, n7482, n7497, n7503, n7510, n7514,
         n7519, n7520, n7524, n7525, n7531, n7538, n7542, n7549, n7552, n7553,
         n7558, n7567, n7574, n7586, n7588, n7603, n7604, n7606, n7611, n7615,
         n7621;
  wire   [511:0] images_bus;
  wire   [8:0] distance;
  wire   [8:0] temp_minimum;
  assign temp_new_reference[0] = N3231;
  assign temp_new_reference[1] = N3232;
  assign temp_new_reference[2] = N3233;
  assign temp_new_reference[3] = N3234;
  assign temp_new_reference[4] = N3235;
  assign N6867 = num_images[0];
  assign N11556 = num_images[8];
  assign count_image[5] = \lt_82/A[5] ;
  assign count_image[4] = \lt_82/A[4] ;
  assign reorder_WEB2 = 1'b1;
  assign reorder_WEB1 = 1'b1;

  dfcrn1 \count_image_reg[4]  ( .D(n12737), .CP(clk), .CDN(n627), .QN(n12188)
         );
  dfcrn1 \count_image_reg[5]  ( .D(n12736), .CP(clk), .CDN(n598), .QN(n12187)
         );
  dfprb1 \distance_reg[8]  ( .D(n13272), .CP(clk), .SDN(n658), .Q(distance[8]), 
        .QN(n12092) );
  dfprb1 \distance_reg[7]  ( .D(n13273), .CP(clk), .SDN(n658), .QN(n12090) );
  dfprb1 \distance_reg[6]  ( .D(n13274), .CP(clk), .SDN(n658), .Q(distance[6]), 
        .QN(n12088) );
  dfprb1 \distance_reg[5]  ( .D(n13275), .CP(clk), .SDN(n658), .Q(distance[5]), 
        .QN(n12086) );
  dfprb1 \distance_reg[4]  ( .D(n13276), .CP(clk), .SDN(n658), .Q(distance[4]), 
        .QN(n12084) );
  dfprb1 \distance_reg[3]  ( .D(n13277), .CP(clk), .SDN(n658), .QN(n12082) );
  dfprb1 \distance_reg[2]  ( .D(n13278), .CP(clk), .SDN(n657), .QN(n12080) );
  dfprb1 \distance_reg[1]  ( .D(n13279), .CP(clk), .SDN(n657), .Q(distance[1]), 
        .QN(n12078) );
  dfprb1 \distance_reg[0]  ( .D(n13280), .CP(clk), .SDN(n657), .QN(n12076) );
  dfprb1 \temp_minimum_reg[0]  ( .D(n13271), .CP(clk), .SDN(n657), .Q(
        temp_minimum[0]), .QN(n12075) );
  dfprb1 \temp_minimum_reg[1]  ( .D(n13270), .CP(clk), .SDN(n658), .QN(n12077)
         );
  dfprb1 \temp_minimum_reg[2]  ( .D(n13269), .CP(clk), .SDN(n657), .Q(
        temp_minimum[2]), .QN(n12079) );
  dfprb1 \temp_minimum_reg[3]  ( .D(n13268), .CP(clk), .SDN(n657), .Q(
        temp_minimum[3]), .QN(n12081) );
  dfprb1 \temp_minimum_reg[4]  ( .D(n13267), .CP(clk), .SDN(n657), .QN(n12083)
         );
  dfprb1 \temp_minimum_reg[5]  ( .D(n13266), .CP(clk), .SDN(n657), .QN(n12085)
         );
  dfprb1 \temp_minimum_reg[6]  ( .D(n13265), .CP(clk), .SDN(n657), .QN(n12087)
         );
  dfprb1 \temp_minimum_reg[7]  ( .D(n13264), .CP(clk), .SDN(n657), .Q(
        temp_minimum[7]), .QN(n12089) );
  dfprb1 \temp_minimum_reg[8]  ( .D(n13263), .CP(clk), .SDN(n656), .Q(
        temp_minimum[8]), .QN(n12091) );
  dfprb1 \temp_new_reference_reg[2]  ( .D(n13260), .CP(clk), .SDN(n656), .Q(
        N3233), .QN(n12210) );
  dfprb1 \temp_new_reference_reg[3]  ( .D(n13259), .CP(clk), .SDN(n656), .Q(
        N3234), .QN(n12209) );
  dfprb1 \temp_new_reference_reg[4]  ( .D(n13258), .CP(clk), .SDN(n656), .Q(
        N3235), .QN(n12208) );
  dfprb1 \temp_new_reference_reg[5]  ( .D(n13257), .CP(clk), .SDN(n656), .Q(
        temp_new_reference[5]), .QN(n12207) );
  dfprb1 \temp_new_reference_reg[6]  ( .D(n13256), .CP(clk), .SDN(n657), .Q(
        temp_new_reference[6]), .QN(n12206) );
  dfprb1 \temp_new_reference_reg[7]  ( .D(n13255), .CP(clk), .SDN(n656), .Q(
        temp_new_reference[7]), .QN(n12205) );
  dfprb1 \temp_new_reference_reg[8]  ( .D(n13254), .CP(clk), .SDN(n656), .Q(
        temp_new_reference[8]), .QN(n12204) );
  dfprb1 \temp_new_reference_reg[1]  ( .D(n13261), .CP(clk), .SDN(n656), .Q(
        N3232), .QN(n12211) );
  dfcrn1 \current_image_index_reg[8]  ( .D(n12725), .CP(clk), .CDN(n620), .QN(
        n12184) );
  dfcrn1 \current_image_index_reg[7]  ( .D(n12726), .CP(clk), .CDN(n612), .QN(
        n12183) );
  dfcrn1 \current_image_index_reg[6]  ( .D(n12727), .CP(clk), .CDN(n613), .QN(
        n12182) );
  dfcrn1 \current_image_index_reg[5]  ( .D(n12728), .CP(clk), .CDN(n613), .QN(
        n12181) );
  dfcrn1 \current_image_index_reg[4]  ( .D(n12729), .CP(clk), .CDN(n613), .QN(
        n12180) );
  dfcrn1 \current_image_index_reg[3]  ( .D(n12730), .CP(clk), .CDN(n613), .QN(
        n12179) );
  dfcrn1 \current_image_index_reg[2]  ( .D(n12731), .CP(clk), .CDN(n613), .QN(
        n12178) );
  dfcrn1 \current_image_index_reg[1]  ( .D(n12732), .CP(clk), .CDN(n613), .QN(
        n12177) );
  dfcrn1 \hash_referance_reg[255]  ( .D(n13281), .CP(clk), .CDN(n613), .QN(
        n12213) );
  dfcrn1 \hash_referance_reg[253]  ( .D(n13282), .CP(clk), .CDN(n613), .QN(
        n12215) );
  dfcrn1 \hash_referance_reg[252]  ( .D(n13283), .CP(clk), .CDN(n613), .QN(
        n12216) );
  dfcrn1 \hash_referance_reg[251]  ( .D(n13284), .CP(clk), .CDN(n613), .QN(
        n12217) );
  dfcrn1 \hash_referance_reg[250]  ( .D(n13285), .CP(clk), .CDN(n614), .QN(
        n12218) );
  dfcrn1 \hash_referance_reg[249]  ( .D(n13286), .CP(clk), .CDN(n614), .QN(
        n12219) );
  dfcrn1 \hash_referance_reg[248]  ( .D(n13287), .CP(clk), .CDN(n614), .QN(
        n12220) );
  dfcrn1 \hash_referance_reg[247]  ( .D(n13288), .CP(clk), .CDN(n614), .QN(
        n12221) );
  dfcrn1 \hash_referance_reg[246]  ( .D(n13289), .CP(clk), .CDN(n614), .QN(
        n12222) );
  dfcrn1 \hash_referance_reg[245]  ( .D(n13290), .CP(clk), .CDN(n614), .QN(
        n12223) );
  dfcrn1 \hash_referance_reg[244]  ( .D(n13291), .CP(clk), .CDN(n614), .QN(
        n12224) );
  dfcrn1 \hash_referance_reg[243]  ( .D(n13292), .CP(clk), .CDN(n614), .QN(
        n12225) );
  dfcrn1 \hash_referance_reg[242]  ( .D(n13293), .CP(clk), .CDN(n614), .QN(
        n12226) );
  dfcrn1 \hash_referance_reg[241]  ( .D(n13294), .CP(clk), .CDN(n614), .QN(
        n12227) );
  dfcrn1 \hash_referance_reg[240]  ( .D(n13295), .CP(clk), .CDN(n615), .QN(
        n12228) );
  dfcrn1 \hash_referance_reg[239]  ( .D(n13296), .CP(clk), .CDN(n615), .QN(
        n12229) );
  dfcrn1 \hash_referance_reg[238]  ( .D(n13297), .CP(clk), .CDN(n615), .QN(
        n12230) );
  dfcrn1 \hash_referance_reg[237]  ( .D(n13298), .CP(clk), .CDN(n615), .QN(
        n12231) );
  dfcrn1 \hash_referance_reg[236]  ( .D(n13299), .CP(clk), .CDN(n615), .QN(
        n12232) );
  dfcrn1 \hash_referance_reg[235]  ( .D(n13300), .CP(clk), .CDN(n615), .QN(
        n12233) );
  dfcrn1 \hash_referance_reg[234]  ( .D(n13301), .CP(clk), .CDN(n615), .QN(
        n12234) );
  dfcrn1 \hash_referance_reg[233]  ( .D(n13302), .CP(clk), .CDN(n615), .QN(
        n12235) );
  dfcrn1 \hash_referance_reg[232]  ( .D(n13303), .CP(clk), .CDN(n615), .QN(
        n12236) );
  dfcrn1 \hash_referance_reg[231]  ( .D(n13304), .CP(clk), .CDN(n615), .QN(
        n12237) );
  dfcrn1 \hash_referance_reg[230]  ( .D(n13305), .CP(clk), .CDN(n616), .QN(
        n12238) );
  dfcrn1 \hash_referance_reg[229]  ( .D(n13306), .CP(clk), .CDN(n616), .QN(
        n12239) );
  dfcrn1 \hash_referance_reg[228]  ( .D(n13307), .CP(clk), .CDN(n616), .QN(
        n12240) );
  dfcrn1 \hash_referance_reg[227]  ( .D(n13308), .CP(clk), .CDN(n616), .QN(
        n12241) );
  dfcrn1 \hash_referance_reg[226]  ( .D(n13309), .CP(clk), .CDN(n616), .QN(
        n12242) );
  dfcrn1 \hash_referance_reg[225]  ( .D(n13310), .CP(clk), .CDN(n616), .QN(
        n12243) );
  dfcrn1 \hash_referance_reg[224]  ( .D(n13311), .CP(clk), .CDN(n616), .QN(
        n12244) );
  dfcrn1 \hash_referance_reg[254]  ( .D(n13536), .CP(clk), .CDN(n616), .QN(
        n12214) );
  dfcrn1 \compare_hash_reg[255]  ( .D(n13537), .CP(clk), .CDN(n616), .QN(
        n12469) );
  dfcrn1 \compare_hash_reg[254]  ( .D(n13538), .CP(clk), .CDN(n616), .QN(
        n12470) );
  dfcrn1 \compare_hash_reg[253]  ( .D(n13539), .CP(clk), .CDN(n617), .QN(
        n12471) );
  dfcrn1 \compare_hash_reg[252]  ( .D(n13540), .CP(clk), .CDN(n617), .QN(
        n12472) );
  dfcrn1 \compare_hash_reg[251]  ( .D(n13541), .CP(clk), .CDN(n617), .QN(
        n12473) );
  dfcrn1 \compare_hash_reg[250]  ( .D(n13542), .CP(clk), .CDN(n617), .QN(
        n12474) );
  dfcrn1 \compare_hash_reg[249]  ( .D(n13543), .CP(clk), .CDN(n617), .QN(
        n12475) );
  dfcrn1 \compare_hash_reg[248]  ( .D(n13544), .CP(clk), .CDN(n617), .QN(
        n12476) );
  dfcrn1 \compare_hash_reg[247]  ( .D(n13545), .CP(clk), .CDN(n617), .QN(
        n12477) );
  dfcrn1 \compare_hash_reg[246]  ( .D(n13546), .CP(clk), .CDN(n617), .QN(
        n12478) );
  dfcrn1 \compare_hash_reg[245]  ( .D(n13547), .CP(clk), .CDN(n617), .QN(
        n12479) );
  dfcrn1 \compare_hash_reg[244]  ( .D(n13548), .CP(clk), .CDN(n617), .QN(
        n12480) );
  dfcrn1 \compare_hash_reg[243]  ( .D(n13549), .CP(clk), .CDN(n618), .QN(
        n12481) );
  dfcrn1 \compare_hash_reg[242]  ( .D(n13550), .CP(clk), .CDN(n618), .QN(
        n12482) );
  dfcrn1 \compare_hash_reg[241]  ( .D(n13551), .CP(clk), .CDN(n618), .QN(
        n12483) );
  dfcrn1 \compare_hash_reg[240]  ( .D(n13552), .CP(clk), .CDN(n618), .QN(
        n12484) );
  dfcrn1 \compare_hash_reg[239]  ( .D(n13553), .CP(clk), .CDN(n618), .QN(
        n12485) );
  dfcrn1 \compare_hash_reg[238]  ( .D(n13554), .CP(clk), .CDN(n618), .QN(
        n12486) );
  dfcrn1 \compare_hash_reg[237]  ( .D(n13555), .CP(clk), .CDN(n618), .QN(
        n12487) );
  dfcrn1 \compare_hash_reg[236]  ( .D(n13556), .CP(clk), .CDN(n618), .QN(
        n12488) );
  dfcrn1 \compare_hash_reg[235]  ( .D(n13557), .CP(clk), .CDN(n618), .QN(
        n12489) );
  dfcrn1 \compare_hash_reg[234]  ( .D(n13558), .CP(clk), .CDN(n618), .QN(
        n12490) );
  dfcrn1 \compare_hash_reg[233]  ( .D(n13559), .CP(clk), .CDN(n619), .QN(
        n12491) );
  dfcrn1 \compare_hash_reg[232]  ( .D(n13560), .CP(clk), .CDN(n619), .QN(
        n12492) );
  dfcrn1 \compare_hash_reg[231]  ( .D(n13561), .CP(clk), .CDN(n619), .QN(
        n12493) );
  dfcrn1 \compare_hash_reg[230]  ( .D(n13562), .CP(clk), .CDN(n619), .QN(
        n12494) );
  dfcrn1 \compare_hash_reg[229]  ( .D(n13563), .CP(clk), .CDN(n619), .QN(
        n12495) );
  dfcrn1 \compare_hash_reg[228]  ( .D(n13564), .CP(clk), .CDN(n619), .QN(
        n12496) );
  dfcrn1 \compare_hash_reg[227]  ( .D(n13565), .CP(clk), .CDN(n619), .QN(
        n12497) );
  dfcrn1 \compare_hash_reg[226]  ( .D(n13566), .CP(clk), .CDN(n619), .QN(
        n12498) );
  dfcrn1 \compare_hash_reg[225]  ( .D(n13567), .CP(clk), .CDN(n619), .QN(
        n12499) );
  dfcrn1 \compare_hash_reg[224]  ( .D(n13568), .CP(clk), .CDN(n619), .QN(
        n12500) );
  dfcrn1 \hash_referance_reg[63]  ( .D(n13472), .CP(clk), .CDN(n620), .QN(
        n12405) );
  dfcrn1 \hash_referance_reg[62]  ( .D(n13473), .CP(clk), .CDN(n620), .QN(
        n12406) );
  dfcrn1 \hash_referance_reg[61]  ( .D(n13474), .CP(clk), .CDN(n620), .QN(
        n12407) );
  dfcrn1 \hash_referance_reg[60]  ( .D(n13475), .CP(clk), .CDN(n620), .QN(
        n12408) );
  dfcrn1 \hash_referance_reg[59]  ( .D(n13476), .CP(clk), .CDN(n620), .QN(
        n12409) );
  dfcrn1 \hash_referance_reg[58]  ( .D(n13477), .CP(clk), .CDN(n620), .QN(
        n12410) );
  dfcrn1 \hash_referance_reg[57]  ( .D(n13478), .CP(clk), .CDN(n620), .QN(
        n12411) );
  dfcrn1 \hash_referance_reg[56]  ( .D(n13479), .CP(clk), .CDN(n620), .QN(
        n12412) );
  dfcrn1 \hash_referance_reg[55]  ( .D(n13480), .CP(clk), .CDN(n620), .QN(
        n12413) );
  dfcrn1 \hash_referance_reg[54]  ( .D(n13481), .CP(clk), .CDN(n621), .QN(
        n12414) );
  dfcrn1 \hash_referance_reg[53]  ( .D(n13482), .CP(clk), .CDN(n621), .QN(
        n12415) );
  dfcrn1 \hash_referance_reg[52]  ( .D(n13483), .CP(clk), .CDN(n621), .QN(
        n12416) );
  dfcrn1 \hash_referance_reg[51]  ( .D(n13484), .CP(clk), .CDN(n621), .QN(
        n12417) );
  dfcrn1 \hash_referance_reg[50]  ( .D(n13485), .CP(clk), .CDN(n621), .QN(
        n12418) );
  dfcrn1 \hash_referance_reg[49]  ( .D(n13486), .CP(clk), .CDN(n621), .QN(
        n12419) );
  dfcrn1 \hash_referance_reg[48]  ( .D(n13487), .CP(clk), .CDN(n621), .QN(
        n12420) );
  dfcrn1 \hash_referance_reg[47]  ( .D(n13488), .CP(clk), .CDN(n621), .QN(
        n12421) );
  dfcrn1 \hash_referance_reg[46]  ( .D(n13489), .CP(clk), .CDN(n621), .QN(
        n12422) );
  dfcrn1 \hash_referance_reg[45]  ( .D(n13490), .CP(clk), .CDN(n621), .QN(
        n12423) );
  dfcrn1 \hash_referance_reg[44]  ( .D(n13491), .CP(clk), .CDN(n622), .QN(
        n12424) );
  dfcrn1 \hash_referance_reg[43]  ( .D(n13492), .CP(clk), .CDN(n622), .QN(
        n12425) );
  dfcrn1 \hash_referance_reg[42]  ( .D(n13493), .CP(clk), .CDN(n622), .QN(
        n12426) );
  dfcrn1 \hash_referance_reg[41]  ( .D(n13494), .CP(clk), .CDN(n622), .QN(
        n12427) );
  dfcrn1 \hash_referance_reg[40]  ( .D(n13495), .CP(clk), .CDN(n622), .QN(
        n12428) );
  dfcrn1 \hash_referance_reg[39]  ( .D(n13496), .CP(clk), .CDN(n622), .QN(
        n12429) );
  dfcrn1 \hash_referance_reg[38]  ( .D(n13497), .CP(clk), .CDN(n622), .QN(
        n12430) );
  dfcrn1 \hash_referance_reg[37]  ( .D(n13498), .CP(clk), .CDN(n622), .QN(
        n12431) );
  dfcrn1 \hash_referance_reg[36]  ( .D(n13499), .CP(clk), .CDN(n622), .QN(
        n12432) );
  dfcrn1 \hash_referance_reg[35]  ( .D(n13500), .CP(clk), .CDN(n622), .QN(
        n12433) );
  dfcrn1 \hash_referance_reg[34]  ( .D(n13501), .CP(clk), .CDN(n623), .QN(
        n12434) );
  dfcrn1 \hash_referance_reg[33]  ( .D(n13502), .CP(clk), .CDN(n623), .QN(
        n12435) );
  dfcrn1 \hash_referance_reg[32]  ( .D(n13503), .CP(clk), .CDN(n623), .QN(
        n12436) );
  dfcrn1 \compare_hash_reg[63]  ( .D(n13728), .CP(clk), .CDN(n623), .QN(n12661) );
  dfcrn1 \compare_hash_reg[62]  ( .D(n13729), .CP(clk), .CDN(n623), .QN(n12662) );
  dfcrn1 \compare_hash_reg[61]  ( .D(n13730), .CP(clk), .CDN(n623), .QN(n12663) );
  dfcrn1 \compare_hash_reg[60]  ( .D(n13731), .CP(clk), .CDN(n623), .QN(n12664) );
  dfcrn1 \compare_hash_reg[59]  ( .D(n13732), .CP(clk), .CDN(n623), .QN(n12665) );
  dfcrn1 \compare_hash_reg[58]  ( .D(n13733), .CP(clk), .CDN(n623), .QN(n12666) );
  dfcrn1 \compare_hash_reg[57]  ( .D(n13734), .CP(clk), .CDN(n623), .QN(n12667) );
  dfcrn1 \compare_hash_reg[56]  ( .D(n13735), .CP(clk), .CDN(n624), .QN(n12668) );
  dfcrn1 \compare_hash_reg[55]  ( .D(n13736), .CP(clk), .CDN(n624), .QN(n12669) );
  dfcrn1 \compare_hash_reg[54]  ( .D(n13737), .CP(clk), .CDN(n624), .QN(n12670) );
  dfcrn1 \compare_hash_reg[53]  ( .D(n13738), .CP(clk), .CDN(n624), .QN(n12671) );
  dfcrn1 \compare_hash_reg[52]  ( .D(n13739), .CP(clk), .CDN(n624), .QN(n12672) );
  dfcrn1 \compare_hash_reg[51]  ( .D(n13740), .CP(clk), .CDN(n624), .QN(n12673) );
  dfcrn1 \compare_hash_reg[50]  ( .D(n13741), .CP(clk), .CDN(n624), .QN(n12674) );
  dfcrn1 \compare_hash_reg[49]  ( .D(n13742), .CP(clk), .CDN(n624), .QN(n12675) );
  dfcrn1 \compare_hash_reg[48]  ( .D(n13743), .CP(clk), .CDN(n624), .QN(n12676) );
  dfcrn1 \compare_hash_reg[47]  ( .D(n13744), .CP(clk), .CDN(n624), .QN(n12677) );
  dfcrn1 \compare_hash_reg[46]  ( .D(n13745), .CP(clk), .CDN(n625), .QN(n12678) );
  dfcrn1 \compare_hash_reg[45]  ( .D(n13746), .CP(clk), .CDN(n625), .QN(n12679) );
  dfcrn1 \compare_hash_reg[44]  ( .D(n13747), .CP(clk), .CDN(n625), .QN(n12680) );
  dfcrn1 \compare_hash_reg[43]  ( .D(n13748), .CP(clk), .CDN(n625), .QN(n12681) );
  dfcrn1 \compare_hash_reg[42]  ( .D(n13749), .CP(clk), .CDN(n625), .QN(n12682) );
  dfcrn1 \compare_hash_reg[41]  ( .D(n13750), .CP(clk), .CDN(n625), .QN(n12683) );
  dfcrn1 \compare_hash_reg[40]  ( .D(n13751), .CP(clk), .CDN(n625), .QN(n12684) );
  dfcrn1 \compare_hash_reg[39]  ( .D(n13752), .CP(clk), .CDN(n625), .QN(n12685) );
  dfcrn1 \compare_hash_reg[38]  ( .D(n13753), .CP(clk), .CDN(n625), .QN(n12686) );
  dfcrn1 \compare_hash_reg[37]  ( .D(n13754), .CP(clk), .CDN(n625), .QN(n12687) );
  dfcrn1 \compare_hash_reg[36]  ( .D(n13755), .CP(clk), .CDN(n626), .QN(n12688) );
  dfcrn1 \compare_hash_reg[35]  ( .D(n13756), .CP(clk), .CDN(n626), .QN(n12689) );
  dfcrn1 \compare_hash_reg[34]  ( .D(n13757), .CP(clk), .CDN(n626), .QN(n12690) );
  dfcrn1 \compare_hash_reg[33]  ( .D(n13758), .CP(clk), .CDN(n626), .QN(n12691) );
  dfcrn1 \compare_hash_reg[32]  ( .D(n13759), .CP(clk), .CDN(n626), .QN(n12692) );
  dfcrn1 \hash_referance_reg[31]  ( .D(n13504), .CP(clk), .CDN(n626), .QN(
        n12437) );
  dfcrn1 \hash_referance_reg[30]  ( .D(n13505), .CP(clk), .CDN(n626), .QN(
        n12438) );
  dfcrn1 \hash_referance_reg[29]  ( .D(n13506), .CP(clk), .CDN(n626), .QN(
        n12439) );
  dfcrn1 \hash_referance_reg[28]  ( .D(n13507), .CP(clk), .CDN(n626), .QN(
        n12440) );
  dfcrn1 \hash_referance_reg[27]  ( .D(n13508), .CP(clk), .CDN(n626), .QN(
        n12441) );
  dfcrn1 \hash_referance_reg[26]  ( .D(n13509), .CP(clk), .CDN(n627), .QN(
        n12442) );
  dfcrn1 \hash_referance_reg[25]  ( .D(n13510), .CP(clk), .CDN(n627), .QN(
        n12443) );
  dfcrn1 \hash_referance_reg[24]  ( .D(n13511), .CP(clk), .CDN(n627), .QN(
        n12444) );
  dfcrn1 \hash_referance_reg[23]  ( .D(n13512), .CP(clk), .CDN(n605), .QN(
        n12445) );
  dfcrn1 \hash_referance_reg[22]  ( .D(n13513), .CP(clk), .CDN(n605), .QN(
        n12446) );
  dfcrn1 \hash_referance_reg[21]  ( .D(n13514), .CP(clk), .CDN(n605), .QN(
        n12447) );
  dfcrn1 \hash_referance_reg[20]  ( .D(n13515), .CP(clk), .CDN(n605), .QN(
        n12448) );
  dfcrn1 \hash_referance_reg[19]  ( .D(n13516), .CP(clk), .CDN(n605), .QN(
        n12449) );
  dfcrn1 \hash_referance_reg[18]  ( .D(n13517), .CP(clk), .CDN(n605), .QN(
        n12450) );
  dfcrn1 \hash_referance_reg[17]  ( .D(n13518), .CP(clk), .CDN(n604), .QN(
        n12451) );
  dfcrn1 \hash_referance_reg[16]  ( .D(n13519), .CP(clk), .CDN(n604), .QN(
        n12452) );
  dfcrn1 \hash_referance_reg[15]  ( .D(n13520), .CP(clk), .CDN(n604), .QN(
        n12453) );
  dfcrn1 \hash_referance_reg[14]  ( .D(n13521), .CP(clk), .CDN(n604), .QN(
        n12454) );
  dfcrn1 \hash_referance_reg[13]  ( .D(n13522), .CP(clk), .CDN(n604), .QN(
        n12455) );
  dfcrn1 \hash_referance_reg[12]  ( .D(n13523), .CP(clk), .CDN(n604), .QN(
        n12456) );
  dfcrn1 \hash_referance_reg[11]  ( .D(n13524), .CP(clk), .CDN(n604), .QN(
        n12457) );
  dfcrn1 \hash_referance_reg[10]  ( .D(n13525), .CP(clk), .CDN(n604), .QN(
        n12458) );
  dfcrn1 \hash_referance_reg[9]  ( .D(n13526), .CP(clk), .CDN(n604), .QN(
        n12459) );
  dfcrn1 \hash_referance_reg[8]  ( .D(n13527), .CP(clk), .CDN(n604), .QN(
        n12460) );
  dfcrn1 \hash_referance_reg[7]  ( .D(n13528), .CP(clk), .CDN(n603), .QN(
        n12461) );
  dfcrn1 \hash_referance_reg[6]  ( .D(n13529), .CP(clk), .CDN(n603), .QN(
        n12462) );
  dfcrn1 \hash_referance_reg[5]  ( .D(n13530), .CP(clk), .CDN(n603), .QN(
        n12463) );
  dfcrn1 \hash_referance_reg[4]  ( .D(n13531), .CP(clk), .CDN(n603), .QN(
        n12464) );
  dfcrn1 \hash_referance_reg[3]  ( .D(n13532), .CP(clk), .CDN(n603), .QN(
        n12465) );
  dfcrn1 \hash_referance_reg[2]  ( .D(n13533), .CP(clk), .CDN(n603), .QN(
        n12466) );
  dfcrn1 \hash_referance_reg[1]  ( .D(n13534), .CP(clk), .CDN(n603), .QN(
        n12467) );
  dfcrn1 \hash_referance_reg[0]  ( .D(n13535), .CP(clk), .CDN(n603), .QN(
        n12468) );
  dfcrn1 \compare_hash_reg[31]  ( .D(n13760), .CP(clk), .CDN(n603), .QN(n12693) );
  dfcrn1 \compare_hash_reg[30]  ( .D(n13761), .CP(clk), .CDN(n603), .QN(n12694) );
  dfcrn1 \compare_hash_reg[29]  ( .D(n13762), .CP(clk), .CDN(n602), .QN(n12695) );
  dfcrn1 \compare_hash_reg[28]  ( .D(n13763), .CP(clk), .CDN(n602), .QN(n12696) );
  dfcrn1 \compare_hash_reg[27]  ( .D(n13764), .CP(clk), .CDN(n602), .QN(n12697) );
  dfcrn1 \compare_hash_reg[26]  ( .D(n13765), .CP(clk), .CDN(n602), .QN(n12698) );
  dfcrn1 \compare_hash_reg[25]  ( .D(n13766), .CP(clk), .CDN(n602), .QN(n12699) );
  dfcrn1 \compare_hash_reg[24]  ( .D(n13767), .CP(clk), .CDN(n602), .QN(n12700) );
  dfcrn1 \compare_hash_reg[23]  ( .D(n13768), .CP(clk), .CDN(n602), .QN(n12701) );
  dfcrn1 \compare_hash_reg[22]  ( .D(n13769), .CP(clk), .CDN(n602), .QN(n12702) );
  dfcrn1 \compare_hash_reg[21]  ( .D(n13770), .CP(clk), .CDN(n602), .QN(n12703) );
  dfcrn1 \compare_hash_reg[20]  ( .D(n13771), .CP(clk), .CDN(n602), .QN(n12704) );
  dfcrn1 \compare_hash_reg[19]  ( .D(n13772), .CP(clk), .CDN(n601), .QN(n12705) );
  dfcrn1 \compare_hash_reg[18]  ( .D(n13773), .CP(clk), .CDN(n601), .QN(n12706) );
  dfcrn1 \compare_hash_reg[17]  ( .D(n13774), .CP(clk), .CDN(n601), .QN(n12707) );
  dfcrn1 \compare_hash_reg[16]  ( .D(n13775), .CP(clk), .CDN(n601), .QN(n12708) );
  dfcrn1 \compare_hash_reg[15]  ( .D(n13776), .CP(clk), .CDN(n601), .QN(n12709) );
  dfcrn1 \compare_hash_reg[14]  ( .D(n13777), .CP(clk), .CDN(n601), .QN(n12710) );
  dfcrn1 \compare_hash_reg[13]  ( .D(n13778), .CP(clk), .CDN(n601), .QN(n12711) );
  dfcrn1 \compare_hash_reg[12]  ( .D(n13779), .CP(clk), .CDN(n601), .QN(n12712) );
  dfcrn1 \compare_hash_reg[11]  ( .D(n13780), .CP(clk), .CDN(n601), .QN(n12713) );
  dfcrn1 \compare_hash_reg[10]  ( .D(n13781), .CP(clk), .CDN(n600), .QN(n12714) );
  dfcrn1 \compare_hash_reg[9]  ( .D(n13782), .CP(clk), .CDN(n600), .QN(n12715)
         );
  dfcrn1 \compare_hash_reg[8]  ( .D(n13783), .CP(clk), .CDN(n600), .QN(n12716)
         );
  dfcrn1 \compare_hash_reg[7]  ( .D(n13784), .CP(clk), .CDN(n600), .QN(n12717)
         );
  dfcrn1 \compare_hash_reg[6]  ( .D(n13785), .CP(clk), .CDN(n600), .QN(n12718)
         );
  dfcrn1 \compare_hash_reg[5]  ( .D(n13786), .CP(clk), .CDN(n600), .QN(n12719)
         );
  dfcrn1 \compare_hash_reg[4]  ( .D(n13787), .CP(clk), .CDN(n600), .QN(n12720)
         );
  dfcrn1 \compare_hash_reg[3]  ( .D(n13788), .CP(clk), .CDN(n600), .QN(n12721)
         );
  dfcrn1 \compare_hash_reg[2]  ( .D(n13789), .CP(clk), .CDN(n600), .QN(n12722)
         );
  dfcrn1 \compare_hash_reg[1]  ( .D(n13790), .CP(clk), .CDN(n600), .QN(n12723)
         );
  dfcrn1 \compare_hash_reg[0]  ( .D(n13791), .CP(clk), .CDN(n599), .QN(n12724)
         );
  dfcrn1 \hash_referance_reg[159]  ( .D(n13376), .CP(clk), .CDN(n599), .QN(
        n12309) );
  dfcrn1 \hash_referance_reg[158]  ( .D(n13377), .CP(clk), .CDN(n599), .QN(
        n12310) );
  dfcrn1 \hash_referance_reg[157]  ( .D(n13378), .CP(clk), .CDN(n599), .QN(
        n12311) );
  dfcrn1 \hash_referance_reg[156]  ( .D(n13379), .CP(clk), .CDN(n599), .QN(
        n12312) );
  dfcrn1 \hash_referance_reg[155]  ( .D(n13380), .CP(clk), .CDN(n599), .QN(
        n12313) );
  dfcrn1 \hash_referance_reg[154]  ( .D(n13381), .CP(clk), .CDN(n599), .QN(
        n12314) );
  dfcrn1 \hash_referance_reg[153]  ( .D(n13382), .CP(clk), .CDN(n599), .QN(
        n12315) );
  dfcrn1 \hash_referance_reg[152]  ( .D(n13383), .CP(clk), .CDN(n599), .QN(
        n12316) );
  dfcrn1 \hash_referance_reg[151]  ( .D(n13384), .CP(clk), .CDN(n599), .QN(
        n12317) );
  dfcrn1 \hash_referance_reg[150]  ( .D(n13385), .CP(clk), .CDN(n598), .QN(
        n12318) );
  dfcrn1 \hash_referance_reg[149]  ( .D(n13386), .CP(clk), .CDN(n598), .QN(
        n12319) );
  dfcrn1 \hash_referance_reg[148]  ( .D(n13387), .CP(clk), .CDN(n598), .QN(
        n12320) );
  dfcrn1 \hash_referance_reg[147]  ( .D(n13388), .CP(clk), .CDN(n598), .QN(
        n12321) );
  dfcrn1 \hash_referance_reg[146]  ( .D(n13389), .CP(clk), .CDN(n598), .QN(
        n12322) );
  dfcrn1 \hash_referance_reg[145]  ( .D(n13390), .CP(clk), .CDN(n598), .QN(
        n12323) );
  dfcrn1 \hash_referance_reg[144]  ( .D(n13391), .CP(clk), .CDN(n601), .QN(
        n12324) );
  dfcrn1 \hash_referance_reg[143]  ( .D(n13392), .CP(clk), .CDN(n605), .QN(
        n12325) );
  dfcrn1 \hash_referance_reg[142]  ( .D(n13393), .CP(clk), .CDN(n605), .QN(
        n12326) );
  dfcrn1 \hash_referance_reg[141]  ( .D(n13394), .CP(clk), .CDN(n605), .QN(
        n12327) );
  dfcrn1 \hash_referance_reg[140]  ( .D(n13395), .CP(clk), .CDN(n605), .QN(
        n12328) );
  dfcrn1 \hash_referance_reg[139]  ( .D(n13396), .CP(clk), .CDN(n606), .QN(
        n12329) );
  dfcrn1 \hash_referance_reg[138]  ( .D(n13397), .CP(clk), .CDN(n606), .QN(
        n12330) );
  dfcrn1 \hash_referance_reg[137]  ( .D(n13398), .CP(clk), .CDN(n606), .QN(
        n12331) );
  dfcrn1 \hash_referance_reg[136]  ( .D(n13399), .CP(clk), .CDN(n606), .QN(
        n12332) );
  dfcrn1 \hash_referance_reg[135]  ( .D(n13400), .CP(clk), .CDN(n606), .QN(
        n12333) );
  dfcrn1 \hash_referance_reg[134]  ( .D(n13401), .CP(clk), .CDN(n606), .QN(
        n12334) );
  dfcrn1 \hash_referance_reg[133]  ( .D(n13402), .CP(clk), .CDN(n606), .QN(
        n12335) );
  dfcrn1 \hash_referance_reg[132]  ( .D(n13403), .CP(clk), .CDN(n606), .QN(
        n12336) );
  dfcrn1 \hash_referance_reg[131]  ( .D(n13404), .CP(clk), .CDN(n606), .QN(
        n12337) );
  dfcrn1 \hash_referance_reg[130]  ( .D(n13405), .CP(clk), .CDN(n606), .QN(
        n12338) );
  dfcrn1 \hash_referance_reg[129]  ( .D(n13406), .CP(clk), .CDN(n607), .QN(
        n12339) );
  dfcrn1 \hash_referance_reg[128]  ( .D(n13407), .CP(clk), .CDN(n607), .QN(
        n12340) );
  dfcrn1 \compare_hash_reg[159]  ( .D(n13632), .CP(clk), .CDN(n607), .QN(
        n12565) );
  dfcrn1 \compare_hash_reg[158]  ( .D(n13633), .CP(clk), .CDN(n607), .QN(
        n12566) );
  dfcrn1 \compare_hash_reg[157]  ( .D(n13634), .CP(clk), .CDN(n607), .QN(
        n12567) );
  dfcrn1 \compare_hash_reg[156]  ( .D(n13635), .CP(clk), .CDN(n607), .QN(
        n12568) );
  dfcrn1 \compare_hash_reg[155]  ( .D(n13636), .CP(clk), .CDN(n607), .QN(
        n12569) );
  dfcrn1 \compare_hash_reg[154]  ( .D(n13637), .CP(clk), .CDN(n607), .QN(
        n12570) );
  dfcrn1 \compare_hash_reg[153]  ( .D(n13638), .CP(clk), .CDN(n607), .QN(
        n12571) );
  dfcrn1 \compare_hash_reg[152]  ( .D(n13639), .CP(clk), .CDN(n607), .QN(
        n12572) );
  dfcrn1 \compare_hash_reg[151]  ( .D(n13640), .CP(clk), .CDN(n608), .QN(
        n12573) );
  dfcrn1 \compare_hash_reg[150]  ( .D(n13641), .CP(clk), .CDN(n608), .QN(
        n12574) );
  dfcrn1 \compare_hash_reg[149]  ( .D(n13642), .CP(clk), .CDN(n608), .QN(
        n12575) );
  dfcrn1 \compare_hash_reg[148]  ( .D(n13643), .CP(clk), .CDN(n608), .QN(
        n12576) );
  dfcrn1 \compare_hash_reg[147]  ( .D(n13644), .CP(clk), .CDN(n608), .QN(
        n12577) );
  dfcrn1 \compare_hash_reg[146]  ( .D(n13645), .CP(clk), .CDN(n608), .QN(
        n12578) );
  dfcrn1 \compare_hash_reg[145]  ( .D(n13646), .CP(clk), .CDN(n608), .QN(
        n12579) );
  dfcrn1 \compare_hash_reg[144]  ( .D(n13647), .CP(clk), .CDN(n608), .QN(
        n12580) );
  dfcrn1 \compare_hash_reg[143]  ( .D(n13648), .CP(clk), .CDN(n608), .QN(
        n12581) );
  dfcrn1 \compare_hash_reg[142]  ( .D(n13649), .CP(clk), .CDN(n608), .QN(
        n12582) );
  dfcrn1 \compare_hash_reg[141]  ( .D(n13650), .CP(clk), .CDN(n609), .QN(
        n12583) );
  dfcrn1 \compare_hash_reg[140]  ( .D(n13651), .CP(clk), .CDN(n609), .QN(
        n12584) );
  dfcrn1 \compare_hash_reg[139]  ( .D(n13652), .CP(clk), .CDN(n609), .QN(
        n12585) );
  dfcrn1 \compare_hash_reg[138]  ( .D(n13653), .CP(clk), .CDN(n609), .QN(
        n12586) );
  dfcrn1 \compare_hash_reg[137]  ( .D(n13654), .CP(clk), .CDN(n609), .QN(
        n12587) );
  dfcrn1 \compare_hash_reg[136]  ( .D(n13655), .CP(clk), .CDN(n609), .QN(
        n12588) );
  dfcrn1 \compare_hash_reg[135]  ( .D(n13656), .CP(clk), .CDN(n609), .QN(
        n12589) );
  dfcrn1 \compare_hash_reg[134]  ( .D(n13657), .CP(clk), .CDN(n609), .QN(
        n12590) );
  dfcrn1 \compare_hash_reg[133]  ( .D(n13658), .CP(clk), .CDN(n609), .QN(
        n12591) );
  dfcrn1 \compare_hash_reg[132]  ( .D(n13659), .CP(clk), .CDN(n609), .QN(
        n12592) );
  dfcrn1 \compare_hash_reg[131]  ( .D(n13660), .CP(clk), .CDN(n610), .QN(
        n12593) );
  dfcrn1 \compare_hash_reg[130]  ( .D(n13661), .CP(clk), .CDN(n610), .QN(
        n12594) );
  dfcrn1 \compare_hash_reg[129]  ( .D(n13662), .CP(clk), .CDN(n610), .QN(
        n12595) );
  dfcrn1 \compare_hash_reg[128]  ( .D(n13663), .CP(clk), .CDN(n610), .QN(
        n12596) );
  dfcrn1 \hash_referance_reg[127]  ( .D(n13408), .CP(clk), .CDN(n610), .QN(
        n12341) );
  dfcrn1 \hash_referance_reg[126]  ( .D(n13409), .CP(clk), .CDN(n610), .QN(
        n12342) );
  dfcrn1 \hash_referance_reg[125]  ( .D(n13410), .CP(clk), .CDN(n610), .QN(
        n12343) );
  dfcrn1 \hash_referance_reg[124]  ( .D(n13411), .CP(clk), .CDN(n610), .QN(
        n12344) );
  dfcrn1 \hash_referance_reg[123]  ( .D(n13412), .CP(clk), .CDN(n610), .QN(
        n12345) );
  dfcrn1 \hash_referance_reg[122]  ( .D(n13413), .CP(clk), .CDN(n610), .QN(
        n12346) );
  dfcrn1 \hash_referance_reg[121]  ( .D(n13414), .CP(clk), .CDN(n611), .QN(
        n12347) );
  dfcrn1 \hash_referance_reg[120]  ( .D(n13415), .CP(clk), .CDN(n611), .QN(
        n12348) );
  dfcrn1 \hash_referance_reg[119]  ( .D(n13416), .CP(clk), .CDN(n611), .QN(
        n12349) );
  dfcrn1 \hash_referance_reg[118]  ( .D(n13417), .CP(clk), .CDN(n611), .QN(
        n12350) );
  dfcrn1 \hash_referance_reg[117]  ( .D(n13418), .CP(clk), .CDN(n611), .QN(
        n12351) );
  dfcrn1 \hash_referance_reg[116]  ( .D(n13419), .CP(clk), .CDN(n611), .QN(
        n12352) );
  dfcrn1 \hash_referance_reg[115]  ( .D(n13420), .CP(clk), .CDN(n611), .QN(
        n12353) );
  dfcrn1 \hash_referance_reg[114]  ( .D(n13421), .CP(clk), .CDN(n611), .QN(
        n12354) );
  dfcrn1 \hash_referance_reg[113]  ( .D(n13422), .CP(clk), .CDN(n611), .QN(
        n12355) );
  dfcrn1 \hash_referance_reg[112]  ( .D(n13423), .CP(clk), .CDN(n611), .QN(
        n12356) );
  dfcrn1 \hash_referance_reg[111]  ( .D(n13424), .CP(clk), .CDN(n612), .QN(
        n12357) );
  dfcrn1 \hash_referance_reg[110]  ( .D(n13425), .CP(clk), .CDN(n612), .QN(
        n12358) );
  dfcrn1 \hash_referance_reg[109]  ( .D(n13426), .CP(clk), .CDN(n612), .QN(
        n12359) );
  dfcrn1 \hash_referance_reg[108]  ( .D(n13427), .CP(clk), .CDN(n612), .QN(
        n12360) );
  dfcrn1 \hash_referance_reg[107]  ( .D(n13428), .CP(clk), .CDN(n612), .QN(
        n12361) );
  dfcrn1 \hash_referance_reg[106]  ( .D(n13429), .CP(clk), .CDN(n612), .QN(
        n12362) );
  dfcrn1 \hash_referance_reg[105]  ( .D(n13430), .CP(clk), .CDN(n612), .QN(
        n12363) );
  dfcrn1 \hash_referance_reg[104]  ( .D(n13431), .CP(clk), .CDN(n612), .QN(
        n12364) );
  dfcrn1 \hash_referance_reg[103]  ( .D(n13432), .CP(clk), .CDN(n612), .QN(
        n12365) );
  dfcrn1 \hash_referance_reg[102]  ( .D(n13433), .CP(clk), .CDN(n652), .QN(
        n12366) );
  dfcrn1 \hash_referance_reg[101]  ( .D(n13434), .CP(clk), .CDN(n641), .QN(
        n12367) );
  dfcrn1 \hash_referance_reg[100]  ( .D(n13435), .CP(clk), .CDN(n641), .QN(
        n12368) );
  dfcrn1 \hash_referance_reg[99]  ( .D(n13436), .CP(clk), .CDN(n642), .QN(
        n12369) );
  dfcrn1 \hash_referance_reg[98]  ( .D(n13437), .CP(clk), .CDN(n642), .QN(
        n12370) );
  dfcrn1 \hash_referance_reg[97]  ( .D(n13438), .CP(clk), .CDN(n642), .QN(
        n12371) );
  dfcrn1 \hash_referance_reg[96]  ( .D(n13439), .CP(clk), .CDN(n642), .QN(
        n12372) );
  dfcrn1 \hash_referance_reg[95]  ( .D(n13440), .CP(clk), .CDN(n642), .QN(
        n12373) );
  dfcrn1 \hash_referance_reg[94]  ( .D(n13441), .CP(clk), .CDN(n642), .QN(
        n12374) );
  dfcrn1 \hash_referance_reg[93]  ( .D(n13442), .CP(clk), .CDN(n642), .QN(
        n12375) );
  dfcrn1 \hash_referance_reg[92]  ( .D(n13443), .CP(clk), .CDN(n642), .QN(
        n12376) );
  dfcrn1 \hash_referance_reg[91]  ( .D(n13444), .CP(clk), .CDN(n642), .QN(
        n12377) );
  dfcrn1 \hash_referance_reg[90]  ( .D(n13445), .CP(clk), .CDN(n642), .QN(
        n12378) );
  dfcrn1 \hash_referance_reg[89]  ( .D(n13446), .CP(clk), .CDN(n643), .QN(
        n12379) );
  dfcrn1 \hash_referance_reg[88]  ( .D(n13447), .CP(clk), .CDN(n643), .QN(
        n12380) );
  dfcrn1 \hash_referance_reg[87]  ( .D(n13448), .CP(clk), .CDN(n643), .QN(
        n12381) );
  dfcrn1 \hash_referance_reg[86]  ( .D(n13449), .CP(clk), .CDN(n643), .QN(
        n12382) );
  dfcrn1 \hash_referance_reg[85]  ( .D(n13450), .CP(clk), .CDN(n643), .QN(
        n12383) );
  dfcrn1 \hash_referance_reg[84]  ( .D(n13451), .CP(clk), .CDN(n643), .QN(
        n12384) );
  dfcrn1 \hash_referance_reg[83]  ( .D(n13452), .CP(clk), .CDN(n643), .QN(
        n12385) );
  dfcrn1 \hash_referance_reg[82]  ( .D(n13453), .CP(clk), .CDN(n643), .QN(
        n12386) );
  dfcrn1 \hash_referance_reg[81]  ( .D(n13454), .CP(clk), .CDN(n643), .QN(
        n12387) );
  dfcrn1 \hash_referance_reg[80]  ( .D(n13455), .CP(clk), .CDN(n643), .QN(
        n12388) );
  dfcrn1 \hash_referance_reg[79]  ( .D(n13456), .CP(clk), .CDN(n644), .QN(
        n12389) );
  dfcrn1 \hash_referance_reg[78]  ( .D(n13457), .CP(clk), .CDN(n644), .QN(
        n12390) );
  dfcrn1 \hash_referance_reg[77]  ( .D(n13458), .CP(clk), .CDN(n644), .QN(
        n12391) );
  dfcrn1 \hash_referance_reg[76]  ( .D(n13459), .CP(clk), .CDN(n644), .QN(
        n12392) );
  dfcrn1 \hash_referance_reg[75]  ( .D(n13460), .CP(clk), .CDN(n644), .QN(
        n12393) );
  dfcrn1 \hash_referance_reg[74]  ( .D(n13461), .CP(clk), .CDN(n644), .QN(
        n12394) );
  dfcrn1 \hash_referance_reg[73]  ( .D(n13462), .CP(clk), .CDN(n644), .QN(
        n12395) );
  dfcrn1 \hash_referance_reg[72]  ( .D(n13463), .CP(clk), .CDN(n644), .QN(
        n12396) );
  dfcrn1 \hash_referance_reg[71]  ( .D(n13464), .CP(clk), .CDN(n644), .QN(
        n12397) );
  dfcrn1 \hash_referance_reg[70]  ( .D(n13465), .CP(clk), .CDN(n644), .QN(
        n12398) );
  dfcrn1 \hash_referance_reg[69]  ( .D(n13466), .CP(clk), .CDN(n645), .QN(
        n12399) );
  dfcrn1 \hash_referance_reg[68]  ( .D(n13467), .CP(clk), .CDN(n645), .QN(
        n12400) );
  dfcrn1 \hash_referance_reg[67]  ( .D(n13468), .CP(clk), .CDN(n645), .QN(
        n12401) );
  dfcrn1 \hash_referance_reg[66]  ( .D(n13469), .CP(clk), .CDN(n645), .QN(
        n12402) );
  dfcrn1 \hash_referance_reg[65]  ( .D(n13470), .CP(clk), .CDN(n645), .QN(
        n12403) );
  dfcrn1 \hash_referance_reg[64]  ( .D(n13471), .CP(clk), .CDN(n645), .QN(
        n12404) );
  dfcrn1 \compare_hash_reg[127]  ( .D(n13664), .CP(clk), .CDN(n645), .QN(
        n12597) );
  dfcrn1 \compare_hash_reg[126]  ( .D(n13665), .CP(clk), .CDN(n645), .QN(
        n12598) );
  dfcrn1 \compare_hash_reg[125]  ( .D(n13666), .CP(clk), .CDN(n645), .QN(
        n12599) );
  dfcrn1 \compare_hash_reg[124]  ( .D(n13667), .CP(clk), .CDN(n645), .QN(
        n12600) );
  dfcrn1 \compare_hash_reg[123]  ( .D(n13668), .CP(clk), .CDN(n646), .QN(
        n12601) );
  dfcrn1 \compare_hash_reg[122]  ( .D(n13669), .CP(clk), .CDN(n646), .QN(
        n12602) );
  dfcrn1 \compare_hash_reg[121]  ( .D(n13670), .CP(clk), .CDN(n646), .QN(
        n12603) );
  dfcrn1 \compare_hash_reg[120]  ( .D(n13671), .CP(clk), .CDN(n646), .QN(
        n12604) );
  dfcrn1 \compare_hash_reg[119]  ( .D(n13672), .CP(clk), .CDN(n646), .QN(
        n12605) );
  dfcrn1 \compare_hash_reg[118]  ( .D(n13673), .CP(clk), .CDN(n646), .QN(
        n12606) );
  dfcrn1 \compare_hash_reg[117]  ( .D(n13674), .CP(clk), .CDN(n646), .QN(
        n12607) );
  dfcrn1 \compare_hash_reg[116]  ( .D(n13675), .CP(clk), .CDN(n646), .QN(
        n12608) );
  dfcrn1 \compare_hash_reg[115]  ( .D(n13676), .CP(clk), .CDN(n646), .QN(
        n12609) );
  dfcrn1 \compare_hash_reg[114]  ( .D(n13677), .CP(clk), .CDN(n646), .QN(
        n12610) );
  dfcrn1 \compare_hash_reg[113]  ( .D(n13678), .CP(clk), .CDN(n647), .QN(
        n12611) );
  dfcrn1 \compare_hash_reg[112]  ( .D(n13679), .CP(clk), .CDN(n647), .QN(
        n12612) );
  dfcrn1 \compare_hash_reg[111]  ( .D(n13680), .CP(clk), .CDN(n647), .QN(
        n12613) );
  dfcrn1 \compare_hash_reg[110]  ( .D(n13681), .CP(clk), .CDN(n647), .QN(
        n12614) );
  dfcrn1 \compare_hash_reg[109]  ( .D(n13682), .CP(clk), .CDN(n647), .QN(
        n12615) );
  dfcrn1 \compare_hash_reg[108]  ( .D(n13683), .CP(clk), .CDN(n647), .QN(
        n12616) );
  dfcrn1 \compare_hash_reg[107]  ( .D(n13684), .CP(clk), .CDN(n647), .QN(
        n12617) );
  dfcrn1 \compare_hash_reg[106]  ( .D(n13685), .CP(clk), .CDN(n647), .QN(
        n12618) );
  dfcrn1 \compare_hash_reg[105]  ( .D(n13686), .CP(clk), .CDN(n647), .QN(
        n12619) );
  dfcrn1 \compare_hash_reg[104]  ( .D(n13687), .CP(clk), .CDN(n647), .QN(
        n12620) );
  dfcrn1 \compare_hash_reg[103]  ( .D(n13688), .CP(clk), .CDN(n648), .QN(
        n12621) );
  dfcrn1 \compare_hash_reg[102]  ( .D(n13689), .CP(clk), .CDN(n648), .QN(
        n12622) );
  dfcrn1 \compare_hash_reg[101]  ( .D(n13690), .CP(clk), .CDN(n648), .QN(
        n12623) );
  dfcrn1 \compare_hash_reg[100]  ( .D(n13691), .CP(clk), .CDN(n648), .QN(
        n12624) );
  dfcrn1 \compare_hash_reg[99]  ( .D(n13692), .CP(clk), .CDN(n648), .QN(n12625) );
  dfcrn1 \compare_hash_reg[98]  ( .D(n13693), .CP(clk), .CDN(n648), .QN(n12626) );
  dfcrn1 \compare_hash_reg[97]  ( .D(n13694), .CP(clk), .CDN(n648), .QN(n12627) );
  dfcrn1 \compare_hash_reg[96]  ( .D(n13695), .CP(clk), .CDN(n648), .QN(n12628) );
  dfcrn1 \compare_hash_reg[95]  ( .D(n13696), .CP(clk), .CDN(n648), .QN(n12629) );
  dfcrn1 \compare_hash_reg[94]  ( .D(n13697), .CP(clk), .CDN(n656), .QN(n12630) );
  dfcrn1 \compare_hash_reg[93]  ( .D(n13698), .CP(clk), .CDN(n656), .QN(n12631) );
  dfcrn1 \compare_hash_reg[92]  ( .D(n13699), .CP(clk), .CDN(n655), .QN(n12632) );
  dfcrn1 \compare_hash_reg[91]  ( .D(n13700), .CP(clk), .CDN(n655), .QN(n12633) );
  dfcrn1 \compare_hash_reg[90]  ( .D(n13701), .CP(clk), .CDN(n655), .QN(n12634) );
  dfcrn1 \compare_hash_reg[89]  ( .D(n13702), .CP(clk), .CDN(n655), .QN(n12635) );
  dfcrn1 \compare_hash_reg[88]  ( .D(n13703), .CP(clk), .CDN(n655), .QN(n12636) );
  dfcrn1 \compare_hash_reg[87]  ( .D(n13704), .CP(clk), .CDN(n655), .QN(n12637) );
  dfcrn1 \compare_hash_reg[86]  ( .D(n13705), .CP(clk), .CDN(n655), .QN(n12638) );
  dfcrn1 \compare_hash_reg[85]  ( .D(n13706), .CP(clk), .CDN(n655), .QN(n12639) );
  dfcrn1 \compare_hash_reg[84]  ( .D(n13707), .CP(clk), .CDN(n655), .QN(n12640) );
  dfcrn1 \compare_hash_reg[83]  ( .D(n13708), .CP(clk), .CDN(n655), .QN(n12641) );
  dfcrn1 \compare_hash_reg[82]  ( .D(n13709), .CP(clk), .CDN(n654), .QN(n12642) );
  dfcrn1 \compare_hash_reg[81]  ( .D(n13710), .CP(clk), .CDN(n654), .QN(n12643) );
  dfcrn1 \compare_hash_reg[80]  ( .D(n13711), .CP(clk), .CDN(n654), .QN(n12644) );
  dfcrn1 \compare_hash_reg[79]  ( .D(n13712), .CP(clk), .CDN(n654), .QN(n12645) );
  dfcrn1 \compare_hash_reg[78]  ( .D(n13713), .CP(clk), .CDN(n654), .QN(n12646) );
  dfcrn1 \compare_hash_reg[77]  ( .D(n13714), .CP(clk), .CDN(n654), .QN(n12647) );
  dfcrn1 \compare_hash_reg[76]  ( .D(n13715), .CP(clk), .CDN(n654), .QN(n12648) );
  dfcrn1 \compare_hash_reg[75]  ( .D(n13716), .CP(clk), .CDN(n654), .QN(n12649) );
  dfcrn1 \compare_hash_reg[74]  ( .D(n13717), .CP(clk), .CDN(n654), .QN(n12650) );
  dfcrn1 \compare_hash_reg[73]  ( .D(n13718), .CP(clk), .CDN(n654), .QN(n12651) );
  dfcrn1 \compare_hash_reg[72]  ( .D(n13719), .CP(clk), .CDN(n653), .QN(n12652) );
  dfcrn1 \compare_hash_reg[71]  ( .D(n13720), .CP(clk), .CDN(n653), .QN(n12653) );
  dfcrn1 \compare_hash_reg[70]  ( .D(n13721), .CP(clk), .CDN(n653), .QN(n12654) );
  dfcrn1 \compare_hash_reg[69]  ( .D(n13722), .CP(clk), .CDN(n653), .QN(n12655) );
  dfcrn1 \compare_hash_reg[68]  ( .D(n13723), .CP(clk), .CDN(n653), .QN(n12656) );
  dfcrn1 \compare_hash_reg[67]  ( .D(n13724), .CP(clk), .CDN(n653), .QN(n12657) );
  dfcrn1 \compare_hash_reg[66]  ( .D(n13725), .CP(clk), .CDN(n653), .QN(n12658) );
  dfcrn1 \compare_hash_reg[65]  ( .D(n13726), .CP(clk), .CDN(n653), .QN(n12659) );
  dfcrn1 \compare_hash_reg[64]  ( .D(n13727), .CP(clk), .CDN(n653), .QN(n12660) );
  dfcrn1 \hash_referance_reg[223]  ( .D(n13312), .CP(clk), .CDN(n653), .QN(
        n12245) );
  dfcrn1 \hash_referance_reg[222]  ( .D(n13313), .CP(clk), .CDN(n652), .QN(
        n12246) );
  dfcrn1 \hash_referance_reg[221]  ( .D(n13314), .CP(clk), .CDN(n652), .QN(
        n12247) );
  dfcrn1 \hash_referance_reg[220]  ( .D(n13315), .CP(clk), .CDN(n652), .QN(
        n12248) );
  dfcrn1 \hash_referance_reg[219]  ( .D(n13316), .CP(clk), .CDN(n652), .QN(
        n12249) );
  dfcrn1 \hash_referance_reg[218]  ( .D(n13317), .CP(clk), .CDN(n652), .QN(
        n12250) );
  dfcrn1 \hash_referance_reg[217]  ( .D(n13318), .CP(clk), .CDN(n652), .QN(
        n12251) );
  dfcrn1 \hash_referance_reg[216]  ( .D(n13319), .CP(clk), .CDN(n652), .QN(
        n12252) );
  dfcrn1 \hash_referance_reg[215]  ( .D(n13320), .CP(clk), .CDN(n652), .QN(
        n12253) );
  dfcrn1 \hash_referance_reg[214]  ( .D(n13321), .CP(clk), .CDN(n652), .QN(
        n12254) );
  dfcrn1 \hash_referance_reg[213]  ( .D(n13322), .CP(clk), .CDN(n651), .QN(
        n12255) );
  dfcrn1 \hash_referance_reg[212]  ( .D(n13323), .CP(clk), .CDN(n651), .QN(
        n12256) );
  dfcrn1 \hash_referance_reg[211]  ( .D(n13324), .CP(clk), .CDN(n651), .QN(
        n12257) );
  dfcrn1 \hash_referance_reg[210]  ( .D(n13325), .CP(clk), .CDN(n651), .QN(
        n12258) );
  dfcrn1 \hash_referance_reg[209]  ( .D(n13326), .CP(clk), .CDN(n651), .QN(
        n12259) );
  dfcrn1 \hash_referance_reg[208]  ( .D(n13327), .CP(clk), .CDN(n651), .QN(
        n12260) );
  dfcrn1 \hash_referance_reg[207]  ( .D(n13328), .CP(clk), .CDN(n651), .QN(
        n12261) );
  dfcrn1 \hash_referance_reg[206]  ( .D(n13329), .CP(clk), .CDN(n651), .QN(
        n12262) );
  dfcrn1 \hash_referance_reg[205]  ( .D(n13330), .CP(clk), .CDN(n651), .QN(
        n12263) );
  dfcrn1 \hash_referance_reg[204]  ( .D(n13331), .CP(clk), .CDN(n651), .QN(
        n12264) );
  dfcrn1 \hash_referance_reg[203]  ( .D(n13332), .CP(clk), .CDN(n650), .QN(
        n12265) );
  dfcrn1 \hash_referance_reg[202]  ( .D(n13333), .CP(clk), .CDN(n650), .QN(
        n12266) );
  dfcrn1 \hash_referance_reg[201]  ( .D(n13334), .CP(clk), .CDN(n650), .QN(
        n12267) );
  dfcrn1 \hash_referance_reg[200]  ( .D(n13335), .CP(clk), .CDN(n650), .QN(
        n12268) );
  dfcrn1 \hash_referance_reg[199]  ( .D(n13336), .CP(clk), .CDN(n650), .QN(
        n12269) );
  dfcrn1 \hash_referance_reg[198]  ( .D(n13337), .CP(clk), .CDN(n650), .QN(
        n12270) );
  dfcrn1 \hash_referance_reg[197]  ( .D(n13338), .CP(clk), .CDN(n650), .QN(
        n12271) );
  dfcrn1 \hash_referance_reg[196]  ( .D(n13339), .CP(clk), .CDN(n650), .QN(
        n12272) );
  dfcrn1 \hash_referance_reg[195]  ( .D(n13340), .CP(clk), .CDN(n650), .QN(
        n12273) );
  dfcrn1 \hash_referance_reg[194]  ( .D(n13341), .CP(clk), .CDN(n650), .QN(
        n12274) );
  dfcrn1 \hash_referance_reg[193]  ( .D(n13342), .CP(clk), .CDN(n649), .QN(
        n12275) );
  dfcrn1 \hash_referance_reg[192]  ( .D(n13343), .CP(clk), .CDN(n649), .QN(
        n12276) );
  dfcrn1 \hash_referance_reg[191]  ( .D(n13344), .CP(clk), .CDN(n649), .QN(
        n12277) );
  dfcrn1 \hash_referance_reg[190]  ( .D(n13345), .CP(clk), .CDN(n649), .QN(
        n12278) );
  dfcrn1 \hash_referance_reg[189]  ( .D(n13346), .CP(clk), .CDN(n649), .QN(
        n12279) );
  dfcrn1 \hash_referance_reg[188]  ( .D(n13347), .CP(clk), .CDN(n649), .QN(
        n12280) );
  dfcrn1 \hash_referance_reg[187]  ( .D(n13348), .CP(clk), .CDN(n649), .QN(
        n12281) );
  dfcrn1 \hash_referance_reg[186]  ( .D(n13349), .CP(clk), .CDN(n649), .QN(
        n12282) );
  dfcrn1 \hash_referance_reg[185]  ( .D(n13350), .CP(clk), .CDN(n649), .QN(
        n12283) );
  dfcrn1 \hash_referance_reg[184]  ( .D(n13351), .CP(clk), .CDN(n649), .QN(
        n12284) );
  dfcrn1 \hash_referance_reg[183]  ( .D(n13352), .CP(clk), .CDN(n648), .QN(
        n12285) );
  dfcrn1 \hash_referance_reg[182]  ( .D(n13353), .CP(clk), .CDN(n634), .QN(
        n12286) );
  dfcrn1 \hash_referance_reg[181]  ( .D(n13354), .CP(clk), .CDN(n627), .QN(
        n12287) );
  dfcrn1 \hash_referance_reg[180]  ( .D(n13355), .CP(clk), .CDN(n627), .QN(
        n12288) );
  dfcrn1 \hash_referance_reg[179]  ( .D(n13356), .CP(clk), .CDN(n627), .QN(
        n12289) );
  dfcrn1 \hash_referance_reg[178]  ( .D(n13357), .CP(clk), .CDN(n627), .QN(
        n12290) );
  dfcrn1 \hash_referance_reg[177]  ( .D(n13358), .CP(clk), .CDN(n627), .QN(
        n12291) );
  dfcrn1 \hash_referance_reg[176]  ( .D(n13359), .CP(clk), .CDN(n627), .QN(
        n12292) );
  dfcrn1 \hash_referance_reg[175]  ( .D(n13360), .CP(clk), .CDN(n628), .QN(
        n12293) );
  dfcrn1 \hash_referance_reg[174]  ( .D(n13361), .CP(clk), .CDN(n628), .QN(
        n12294) );
  dfcrn1 \hash_referance_reg[173]  ( .D(n13362), .CP(clk), .CDN(n628), .QN(
        n12295) );
  dfcrn1 \hash_referance_reg[172]  ( .D(n13363), .CP(clk), .CDN(n628), .QN(
        n12296) );
  dfcrn1 \hash_referance_reg[171]  ( .D(n13364), .CP(clk), .CDN(n628), .QN(
        n12297) );
  dfcrn1 \hash_referance_reg[170]  ( .D(n13365), .CP(clk), .CDN(n628), .QN(
        n12298) );
  dfcrn1 \hash_referance_reg[169]  ( .D(n13366), .CP(clk), .CDN(n628), .QN(
        n12299) );
  dfcrn1 \hash_referance_reg[168]  ( .D(n13367), .CP(clk), .CDN(n628), .QN(
        n12300) );
  dfcrn1 \hash_referance_reg[167]  ( .D(n13368), .CP(clk), .CDN(n628), .QN(
        n12301) );
  dfcrn1 \hash_referance_reg[166]  ( .D(n13369), .CP(clk), .CDN(n628), .QN(
        n12302) );
  dfcrn1 \hash_referance_reg[165]  ( .D(n13370), .CP(clk), .CDN(n629), .QN(
        n12303) );
  dfcrn1 \hash_referance_reg[164]  ( .D(n13371), .CP(clk), .CDN(n629), .QN(
        n12304) );
  dfcrn1 \hash_referance_reg[163]  ( .D(n13372), .CP(clk), .CDN(n629), .QN(
        n12305) );
  dfcrn1 \hash_referance_reg[162]  ( .D(n13373), .CP(clk), .CDN(n629), .QN(
        n12306) );
  dfcrn1 \hash_referance_reg[161]  ( .D(n13374), .CP(clk), .CDN(n629), .QN(
        n12307) );
  dfcrn1 \hash_referance_reg[160]  ( .D(n13375), .CP(clk), .CDN(n629), .QN(
        n12308) );
  dfcrn1 \compare_hash_reg[223]  ( .D(n13569), .CP(clk), .CDN(n629), .QN(
        n12501) );
  dfcrn1 \compare_hash_reg[222]  ( .D(n13570), .CP(clk), .CDN(n629), .QN(
        n12502) );
  dfcrn1 \compare_hash_reg[221]  ( .D(n13571), .CP(clk), .CDN(n629), .QN(
        n12503) );
  dfcrn1 \compare_hash_reg[220]  ( .D(n13572), .CP(clk), .CDN(n629), .QN(
        n12504) );
  dfcrn1 \compare_hash_reg[219]  ( .D(n13573), .CP(clk), .CDN(n630), .QN(
        n12505) );
  dfcrn1 \compare_hash_reg[218]  ( .D(n13574), .CP(clk), .CDN(n630), .QN(
        n12506) );
  dfcrn1 \compare_hash_reg[217]  ( .D(n13575), .CP(clk), .CDN(n630), .QN(
        n12507) );
  dfcrn1 \compare_hash_reg[216]  ( .D(n13576), .CP(clk), .CDN(n630), .QN(
        n12508) );
  dfcrn1 \compare_hash_reg[215]  ( .D(n13577), .CP(clk), .CDN(n630), .QN(
        n12509) );
  dfcrn1 \compare_hash_reg[214]  ( .D(n13578), .CP(clk), .CDN(n630), .QN(
        n12510) );
  dfcrn1 \compare_hash_reg[213]  ( .D(n13579), .CP(clk), .CDN(n630), .QN(
        n12511) );
  dfcrn1 \compare_hash_reg[212]  ( .D(n13580), .CP(clk), .CDN(n630), .QN(
        n12512) );
  dfcrn1 \compare_hash_reg[211]  ( .D(n13581), .CP(clk), .CDN(n630), .QN(
        n12513) );
  dfcrn1 \compare_hash_reg[210]  ( .D(n13582), .CP(clk), .CDN(n630), .QN(
        n12514) );
  dfcrn1 \compare_hash_reg[209]  ( .D(n13583), .CP(clk), .CDN(n631), .QN(
        n12515) );
  dfcrn1 \compare_hash_reg[208]  ( .D(n13584), .CP(clk), .CDN(n631), .QN(
        n12516) );
  dfcrn1 \compare_hash_reg[207]  ( .D(n13585), .CP(clk), .CDN(n631), .QN(
        n12517) );
  dfcrn1 \compare_hash_reg[206]  ( .D(n13586), .CP(clk), .CDN(n631), .QN(
        n12518) );
  dfcrn1 \compare_hash_reg[205]  ( .D(n13587), .CP(clk), .CDN(n631), .QN(
        n12519) );
  dfcrn1 \compare_hash_reg[204]  ( .D(n13588), .CP(clk), .CDN(n631), .QN(
        n12520) );
  dfcrn1 \compare_hash_reg[203]  ( .D(n13589), .CP(clk), .CDN(n631), .QN(
        n12521) );
  dfcrn1 \compare_hash_reg[202]  ( .D(n13590), .CP(clk), .CDN(n631), .QN(
        n12522) );
  dfcrn1 \compare_hash_reg[201]  ( .D(n13591), .CP(clk), .CDN(n631), .QN(
        n12523) );
  dfcrn1 \compare_hash_reg[200]  ( .D(n13592), .CP(clk), .CDN(n631), .QN(
        n12524) );
  dfcrn1 \compare_hash_reg[199]  ( .D(n13593), .CP(clk), .CDN(n632), .QN(
        n12525) );
  dfcrn1 \compare_hash_reg[198]  ( .D(n13594), .CP(clk), .CDN(n632), .QN(
        n12526) );
  dfcrn1 \compare_hash_reg[197]  ( .D(n13595), .CP(clk), .CDN(n632), .QN(
        n12527) );
  dfcrn1 \compare_hash_reg[195]  ( .D(n13596), .CP(clk), .CDN(n632), .QN(
        n12529) );
  dfcrn1 \compare_hash_reg[194]  ( .D(n13597), .CP(clk), .CDN(n632), .QN(
        n12530) );
  dfcrn1 \compare_hash_reg[193]  ( .D(n13598), .CP(clk), .CDN(n632), .QN(
        n12531) );
  dfcrn1 \compare_hash_reg[192]  ( .D(n13599), .CP(clk), .CDN(n632), .QN(
        n12532) );
  dfcrn1 \compare_hash_reg[191]  ( .D(n13600), .CP(clk), .CDN(n632), .QN(
        n12533) );
  dfcrn1 \compare_hash_reg[190]  ( .D(n13601), .CP(clk), .CDN(n632), .QN(
        n12534) );
  dfcrn1 \compare_hash_reg[189]  ( .D(n13602), .CP(clk), .CDN(n632), .QN(
        n12535) );
  dfcrn1 \compare_hash_reg[188]  ( .D(n13603), .CP(clk), .CDN(n633), .QN(
        n12536) );
  dfcrn1 \compare_hash_reg[187]  ( .D(n13604), .CP(clk), .CDN(n633), .QN(
        n12537) );
  dfcrn1 \compare_hash_reg[186]  ( .D(n13605), .CP(clk), .CDN(n633), .QN(
        n12538) );
  dfcrn1 \compare_hash_reg[185]  ( .D(n13606), .CP(clk), .CDN(n633), .QN(
        n12539) );
  dfcrn1 \compare_hash_reg[184]  ( .D(n13607), .CP(clk), .CDN(n633), .QN(
        n12540) );
  dfcrn1 \compare_hash_reg[183]  ( .D(n13608), .CP(clk), .CDN(n633), .QN(
        n12541) );
  dfcrn1 \compare_hash_reg[182]  ( .D(n13609), .CP(clk), .CDN(n633), .QN(
        n12542) );
  dfcrn1 \compare_hash_reg[181]  ( .D(n13610), .CP(clk), .CDN(n633), .QN(
        n12543) );
  dfcrn1 \compare_hash_reg[180]  ( .D(n13611), .CP(clk), .CDN(n633), .QN(
        n12544) );
  dfcrn1 \compare_hash_reg[179]  ( .D(n13612), .CP(clk), .CDN(n633), .QN(
        n12545) );
  dfcrn1 \compare_hash_reg[178]  ( .D(n13613), .CP(clk), .CDN(n634), .QN(
        n12546) );
  dfcrn1 \compare_hash_reg[177]  ( .D(n13614), .CP(clk), .CDN(n634), .QN(
        n12547) );
  dfcrn1 \compare_hash_reg[176]  ( .D(n13615), .CP(clk), .CDN(n634), .QN(
        n12548) );
  dfcrn1 \compare_hash_reg[175]  ( .D(n13616), .CP(clk), .CDN(n634), .QN(
        n12549) );
  dfcrn1 \compare_hash_reg[174]  ( .D(n13617), .CP(clk), .CDN(n634), .QN(
        n12550) );
  dfcrn1 \compare_hash_reg[173]  ( .D(n13618), .CP(clk), .CDN(n634), .QN(
        n12551) );
  dfcrn1 \compare_hash_reg[172]  ( .D(n13619), .CP(clk), .CDN(n634), .QN(
        n12552) );
  dfcrn1 \compare_hash_reg[171]  ( .D(n13620), .CP(clk), .CDN(n634), .QN(
        n12553) );
  dfcrn1 \compare_hash_reg[170]  ( .D(n13621), .CP(clk), .CDN(n634), .QN(
        n12554) );
  dfcrn1 \compare_hash_reg[169]  ( .D(n13622), .CP(clk), .CDN(n635), .QN(
        n12555) );
  dfcrn1 \compare_hash_reg[168]  ( .D(n13623), .CP(clk), .CDN(n635), .QN(
        n12556) );
  dfcrn1 \compare_hash_reg[167]  ( .D(n13624), .CP(clk), .CDN(n635), .QN(
        n12557) );
  dfcrn1 \compare_hash_reg[166]  ( .D(n13625), .CP(clk), .CDN(n635), .QN(
        n12558) );
  dfcrn1 \compare_hash_reg[165]  ( .D(n13626), .CP(clk), .CDN(n635), .QN(
        n12559) );
  dfcrn1 \compare_hash_reg[164]  ( .D(n13627), .CP(clk), .CDN(n635), .QN(
        n12560) );
  dfcrn1 \compare_hash_reg[163]  ( .D(n13628), .CP(clk), .CDN(n635), .QN(
        n12561) );
  dfcrn1 \compare_hash_reg[162]  ( .D(n13629), .CP(clk), .CDN(n635), .QN(
        n12562) );
  dfcrn1 \compare_hash_reg[161]  ( .D(n13630), .CP(clk), .CDN(n635), .QN(
        n12563) );
  dfcrn1 \compare_hash_reg[160]  ( .D(n13631), .CP(clk), .CDN(n635), .QN(
        n12564) );
  dfcrn1 \compare_hash_reg[196]  ( .D(n13792), .CP(clk), .CDN(n636), .QN(
        n12528) );
  dfprb1 \temp_new_reference_reg[0]  ( .D(n13262), .CP(clk), .SDN(n656), .Q(
        N3231), .QN(n12212) );
  dfcrn1 \current_image_index_reg[0]  ( .D(n12733), .CP(clk), .CDN(n636), .QN(
        n12174) );
  dfcrn1 \images_bus_reg[501]  ( .D(n12752), .CP(clk), .CDN(n636), .QN(n12173)
         );
  dfcrn1 \images_bus_reg[53]  ( .D(n13200), .CP(clk), .CDN(n636), .QN(n12172)
         );
  dfcrn1 \images_bus_reg[397]  ( .D(n12856), .CP(clk), .CDN(n636), .QN(n12171)
         );
  dfcrn1 \images_bus_reg[197]  ( .D(n13056), .CP(clk), .CDN(n636), .QN(n12170)
         );
  dfcrn1 \images_bus_reg[283]  ( .D(n12970), .CP(clk), .CDN(n641), .QN(n12169)
         );
  dfcrn1 \images_bus_reg[187]  ( .D(n13066), .CP(clk), .CDN(n636), .QN(n12168)
         );
  dfcrn1 \images_bus_reg[441]  ( .D(n12812), .CP(clk), .CDN(n636), .QN(n12167)
         );
  dfcrn1 \images_bus_reg[489]  ( .D(n12764), .CP(clk), .CDN(n636), .QN(n12166)
         );
  dfcrn1 \images_bus_reg[361]  ( .D(n12892), .CP(clk), .CDN(n636), .QN(n12165)
         );
  dfcrn1 \images_bus_reg[9]  ( .D(n13244), .CP(clk), .CDN(n637), .QN(n12164)
         );
  dfcrn1 \images_bus_reg[511]  ( .D(n13253), .CP(clk), .CDN(n637), .QN(n12163)
         );
  dfcrn1 \images_bus_reg[510]  ( .D(n12743), .CP(clk), .CDN(n637), .QN(n12162)
         );
  dfcrn1 \images_bus_reg[478]  ( .D(n12775), .CP(clk), .CDN(n637), .QN(n12161)
         );
  dfcrn1 \images_bus_reg[446]  ( .D(n12807), .CP(clk), .CDN(n637), .QN(n12160)
         );
  dfcrn1 \images_bus_reg[190]  ( .D(n13063), .CP(clk), .CDN(n637), .QN(n12159)
         );
  dfcrn1 \images_bus_reg[470]  ( .D(n12783), .CP(clk), .CDN(n637), .QN(n12158)
         );
  dfcrn1 \images_bus_reg[342]  ( .D(n12911), .CP(clk), .CDN(n637), .QN(n12157)
         );
  dfcrn1 \images_bus_reg[462]  ( .D(n12791), .CP(clk), .CDN(n637), .QN(n12156)
         );
  dfcrn1 \images_bus_reg[206]  ( .D(n13047), .CP(clk), .CDN(n637), .QN(n12155)
         );
  dfcrn1 \images_bus_reg[174]  ( .D(n13079), .CP(clk), .CDN(n638), .QN(n12154)
         );
  dfcrn1 \images_bus_reg[294]  ( .D(n12959), .CP(clk), .CDN(n638), .QN(n12153)
         );
  dfcrn1 \images_bus_reg[508]  ( .D(n12745), .CP(clk), .CDN(n638), .QN(n12152)
         );
  dfcrn1 \images_bus_reg[476]  ( .D(n12777), .CP(clk), .CDN(n638), .QN(n12151)
         );
  dfcrn1 \images_bus_reg[412]  ( .D(n12841), .CP(clk), .CDN(n638), .QN(n12150)
         );
  dfcrn1 \images_bus_reg[284]  ( .D(n12969), .CP(clk), .CDN(n638), .QN(n12149)
         );
  dfcrn1 \images_bus_reg[92]  ( .D(n13161), .CP(clk), .CDN(n638), .QN(n12148)
         );
  dfcrn1 \images_bus_reg[468]  ( .D(n12785), .CP(clk), .CDN(n638), .QN(n12147)
         );
  dfcrn1 \images_bus_reg[308]  ( .D(n12945), .CP(clk), .CDN(n638), .QN(n12146)
         );
  dfcrn1 \images_bus_reg[180]  ( .D(n13073), .CP(clk), .CDN(n638), .QN(n12145)
         );
  dfcrn1 \images_bus_reg[148]  ( .D(n13105), .CP(clk), .CDN(n639), .QN(n12144)
         );
  dfcrn1 \images_bus_reg[116]  ( .D(n13137), .CP(clk), .CDN(n639), .QN(n12143)
         );
  dfcrn1 \images_bus_reg[428]  ( .D(n12825), .CP(clk), .CDN(n639), .QN(n12142)
         );
  dfcrn1 \images_bus_reg[452]  ( .D(n12801), .CP(clk), .CDN(n639), .QN(n12141)
         );
  dfcrn1 \images_bus_reg[420]  ( .D(n12833), .CP(clk), .CDN(n639), .QN(n12140)
         );
  dfcrn1 \images_bus_reg[388]  ( .D(n12865), .CP(clk), .CDN(n639), .QN(n12139)
         );
  dfcrn1 \images_bus_reg[356]  ( .D(n12897), .CP(clk), .CDN(n639), .QN(n12138)
         );
  dfcrn1 \images_bus_reg[228]  ( .D(n13025), .CP(clk), .CDN(n639), .QN(n12137)
         );
  dfcrn1 \images_bus_reg[410]  ( .D(n12843), .CP(clk), .CDN(n639), .QN(n12136)
         );
  dfcrn1 \images_bus_reg[378]  ( .D(n12875), .CP(clk), .CDN(n639), .QN(n12135)
         );
  dfcrn1 \images_bus_reg[218]  ( .D(n13035), .CP(clk), .CDN(n640), .QN(n12134)
         );
  dfcrn1 \images_bus_reg[90]  ( .D(n13163), .CP(clk), .CDN(n640), .QN(n12133)
         );
  dfcrn1 \images_bus_reg[370]  ( .D(n12883), .CP(clk), .CDN(n640), .QN(n12132)
         );
  dfcrn1 \images_bus_reg[114]  ( .D(n13139), .CP(clk), .CDN(n640), .QN(n12131)
         );
  dfcrn1 \images_bus_reg[50]  ( .D(n13203), .CP(clk), .CDN(n640), .QN(n12130)
         );
  dfcrn1 \images_bus_reg[458]  ( .D(n12795), .CP(clk), .CDN(n640), .QN(n12129)
         );
  dfcrn1 \images_bus_reg[202]  ( .D(n13051), .CP(clk), .CDN(n640), .QN(n12128)
         );
  dfcrn1 \images_bus_reg[138]  ( .D(n13115), .CP(clk), .CDN(n640), .QN(n12127)
         );
  dfcrn1 \images_bus_reg[10]  ( .D(n13243), .CP(clk), .CDN(n640), .QN(n12126)
         );
  dfcrn1 \images_bus_reg[482]  ( .D(n12771), .CP(clk), .CDN(n640), .QN(n12125)
         );
  dfcrn1 \images_bus_reg[386]  ( .D(n12867), .CP(clk), .CDN(n641), .QN(n12124)
         );
  dfcrn1 \images_bus_reg[354]  ( .D(n12899), .CP(clk), .CDN(n641), .QN(n12123)
         );
  dfcrn1 \images_bus_reg[290]  ( .D(n12963), .CP(clk), .CDN(n641), .QN(n12122)
         );
  dfcrn1 \images_bus_reg[226]  ( .D(n13027), .CP(clk), .CDN(n641), .QN(n12121)
         );
  dfcrn1 \images_bus_reg[34]  ( .D(n13219), .CP(clk), .CDN(n641), .QN(n12120)
         );
  dfcrn1 \images_bus_reg[432]  ( .D(n12821), .CP(clk), .CDN(n641), .QN(n12119)
         );
  dfcrn1 \images_bus_reg[232]  ( .D(n13021), .CP(clk), .CDN(n641), .QN(n12118)
         );
  lanhq1 \last_image_reg[8]  ( .E(N26357), .D(N26366), .Q(last_image[8]) );
  lanhq1 \last_image_reg[7]  ( .E(N26357), .D(N26365), .Q(last_image[7]) );
  lanhq1 \last_image_reg[6]  ( .E(N26357), .D(N26364), .Q(last_image[6]) );
  lanhq1 \last_image_reg[5]  ( .E(N26357), .D(N26363), .Q(last_image[5]) );
  lanhq1 \last_image_reg[4]  ( .E(N26357), .D(N26362), .Q(last_image[4]) );
  lanhq1 \last_image_reg[3]  ( .E(N26357), .D(N26361), .Q(last_image[3]) );
  lanhq1 \last_image_reg[2]  ( .E(N26357), .D(N26360), .Q(last_image[2]) );
  lanhq1 \last_image_reg[1]  ( .E(N26357), .D(N26359), .Q(last_image[1]) );
  lanhq1 \last_image_reg[0]  ( .E(N26357), .D(N26358), .Q(last_image[0]) );
  aon211d1 U7 ( .C1(n3589), .C2(n2754), .B(n3590), .A(reorder_A2[0]), .ZN(
        n3578) );
  aoi222d1 U15 ( .A1(N5070), .A2(n3583), .B1(N3231), .B2(n3593), .C1(N3879), 
        .C2(n951), .ZN(n3598) );
  aoi222d1 U16 ( .A1(reorder_A2[3]), .A2(n3594), .B1(N4688), .B2(n953), .C1(
        N3972), .C2(n1), .ZN(n3597) );
  aoi222d1 U18 ( .A1(N5071), .A2(n3583), .B1(N3232), .B2(n3593), .C1(N3880), 
        .C2(n951), .ZN(n3600) );
  aoi222d1 U19 ( .A1(reorder_A2[4]), .A2(n3594), .B1(N4689), .B2(n952), .C1(
        N3973), .C2(n1), .ZN(n3599) );
  aoi222d1 U1043 ( .A1(N5072), .A2(n3583), .B1(N3233), .B2(n3593), .C1(N3881), 
        .C2(n951), .ZN(n3602) );
  aoi222d1 U1044 ( .A1(reorder_A2[5]), .A2(n3594), .B1(N4690), .B2(n952), .C1(
        n502), .C2(n1), .ZN(n3601) );
  aoi222d1 U1059 ( .A1(N5073), .A2(n3583), .B1(N3234), .B2(n3593), .C1(N3882), 
        .C2(n950), .ZN(n3604) );
  aoi222d1 U1060 ( .A1(reorder_A2[6]), .A2(n3594), .B1(N4691), .B2(n952), .C1(
        n955), .C2(n1), .ZN(n3603) );
  aoi222d1 U1062 ( .A1(N5074), .A2(n3583), .B1(N3235), .B2(n3593), .C1(N3883), 
        .C2(n950), .ZN(n3606) );
  aoi222d1 U1063 ( .A1(reorder_A2[7]), .A2(n3594), .B1(N4692), .B2(n952), .C1(
        N3976), .C2(n1), .ZN(n3605) );
  aoi222d1 U1065 ( .A1(n505), .A2(n1), .B1(N5108), .B2(n3583), .C1(N4693), 
        .C2(n954), .ZN(n3610) );
  oai211d1 U1067 ( .C1(n2783), .C2(n12207), .A(n2754), .B(n3588), .ZN(n3608)
         );
  aon211d1 U1068 ( .C1(n3589), .C2(n2754), .B(n3590), .A(reorder_A2[8]), .ZN(
        n3607) );
  aoi222d1 U1070 ( .A1(N5109), .A2(n3583), .B1(N3237), .B2(n3593), .C1(N3885), 
        .C2(n950), .ZN(n3612) );
  aoi222d1 U1071 ( .A1(reorder_A2[9]), .A2(n3594), .B1(N4694), .B2(n952), .C1(
        N4002), .C2(n1), .ZN(n3611) );
  aoi222d1 U1073 ( .A1(N5110), .A2(n3583), .B1(N3238), .B2(n3593), .C1(N3886), 
        .C2(n950), .ZN(n3614) );
  aoi222d1 U1074 ( .A1(reorder_A2[10]), .A2(n3594), .B1(N4695), .B2(n952), 
        .C1(N4003), .C2(n1), .ZN(n3613) );
  aoi222d1 U1076 ( .A1(N5111), .A2(n3583), .B1(N3239), .B2(n3593), .C1(N3887), 
        .C2(n950), .ZN(n3616) );
  aoi222d1 U1079 ( .A1(reorder_A2[11]), .A2(n3594), .B1(N4696), .B2(n952), 
        .C1(N4004), .C2(n1), .ZN(n3615) );
  aoi222d1 U1091 ( .A1(N5070), .A2(n3583), .B1(N3207), .B2(n3622), .C1(N3843), 
        .C2(n950), .ZN(n3629) );
  aoi222d1 U1092 ( .A1(reorder_A1[3]), .A2(n3623), .B1(N4652), .B2(n952), .C1(
        N3972), .C2(n1), .ZN(n3628) );
  aoi222d1 U1094 ( .A1(N5071), .A2(n3583), .B1(N3208), .B2(n3622), .C1(N3844), 
        .C2(n950), .ZN(n3631) );
  aoi222d1 U1095 ( .A1(reorder_A1[4]), .A2(n3623), .B1(N4653), .B2(n952), .C1(
        N3973), .C2(n1), .ZN(n3630) );
  aoi222d1 U1097 ( .A1(N5072), .A2(n3583), .B1(N3209), .B2(n3622), .C1(N3845), 
        .C2(n950), .ZN(n3633) );
  aoi222d1 U1098 ( .A1(reorder_A1[5]), .A2(n3623), .B1(N4654), .B2(n953), .C1(
        n502), .C2(n1), .ZN(n3632) );
  aoi222d1 U1100 ( .A1(N5073), .A2(n3583), .B1(N3210), .B2(n3622), .C1(N3846), 
        .C2(n950), .ZN(n3635) );
  aoi222d1 U1101 ( .A1(reorder_A1[6]), .A2(n3623), .B1(N4655), .B2(n953), .C1(
        n955), .C2(n1), .ZN(n3634) );
  aoi222d1 U1103 ( .A1(N5074), .A2(n3583), .B1(N3211), .B2(n3622), .C1(N3847), 
        .C2(n950), .ZN(n3637) );
  aoi222d1 U1104 ( .A1(reorder_A1[7]), .A2(n3623), .B1(N4656), .B2(n953), .C1(
        N3976), .C2(n1), .ZN(n3636) );
  aoi222d1 U1106 ( .A1(N5108), .A2(n3583), .B1(N3212), .B2(n3622), .C1(N3848), 
        .C2(n950), .ZN(n3639) );
  aoi222d1 U1107 ( .A1(reorder_A1[8]), .A2(n3623), .B1(N4657), .B2(n953), .C1(
        n505), .C2(n1), .ZN(n3638) );
  aoi222d1 U1109 ( .A1(N5076), .A2(n3583), .B1(N3213), .B2(n3622), .C1(N3849), 
        .C2(n949), .ZN(n3641) );
  aoi222d1 U1110 ( .A1(reorder_A1[9]), .A2(n3623), .B1(N4658), .B2(n953), .C1(
        N3978), .C2(n1), .ZN(n3640) );
  aoi222d1 U1112 ( .A1(N5077), .A2(n3583), .B1(N3214), .B2(n3622), .C1(N3850), 
        .C2(n949), .ZN(n3643) );
  aoi222d1 U1113 ( .A1(reorder_A1[10]), .A2(n3623), .B1(N4659), .B2(n953), 
        .C1(N3979), .C2(n1), .ZN(n3642) );
  aoi222d1 U1115 ( .A1(N5078), .A2(n3583), .B1(N3215), .B2(n3622), .C1(N3851), 
        .C2(n949), .ZN(n3645) );
  aoi222d1 U1121 ( .A1(reorder_A1[11]), .A2(n3623), .B1(N4660), .B2(n953), 
        .C1(N3980), .C2(n1), .ZN(n3644) );
  aor21d1 U1132 ( .B1(n493), .B2(n3657), .A(finish_reordering), .Z(n12117) );
  aor222d1 U1134 ( .A1(N3878), .A2(n3658), .B1(N3914), .B2(n2766), .C1(N4723), 
        .C2(n2), .Z(n12176) );
  oai222d1 U1136 ( .A1(n2780), .A2(n3662), .B1(N3877), .B2(n3663), .C1(n2780), 
        .C2(n2768), .ZN(n3661) );
  aoi31d1 U1137 ( .B1(n2775), .B2(n2777), .B3(n3666), .A(n3667), .ZN(n3663) );
  oai21d1 U1138 ( .B1(reading_current), .B2(reading_compare), .A(n2776), .ZN(
        n3666) );
  oan211d1 U1140 ( .C1(n3670), .C2(n3667), .B(reading_current), .A(n497), .ZN(
        n3669) );
  oai21d1 U1141 ( .B1(n493), .B2(n2782), .A(n3673), .ZN(n12189) );
  aon211d1 U1142 ( .C1(n3674), .C2(N5122), .B(n3657), .A(n493), .ZN(n3673) );
  aoi21d1 U1143 ( .B1(n2774), .B2(n3676), .A(new_reference_is_done), .ZN(n3674) );
  aor22d1 U1144 ( .A1(n500), .A2(n3677), .B1(N5071), .B2(n2755), .Z(n12190) );
  aor22d1 U1145 ( .A1(n502), .A2(n3677), .B1(N5072), .B2(n2755), .Z(n12191) );
  aor22d1 U1146 ( .A1(n955), .A2(n3677), .B1(N5073), .B2(n2755), .Z(n12192) );
  aor22d1 U1147 ( .A1(n504), .A2(n3677), .B1(N5074), .B2(n2755), .Z(n12193) );
  aor22d1 U1148 ( .A1(n506), .A2(n3677), .B1(N4010), .B2(n2755), .Z(n12194) );
  aor22d1 U1149 ( .A1(n508), .A2(n3677), .B1(N4011), .B2(n2755), .Z(n12195) );
  aor22d1 U1150 ( .A1(n509), .A2(n3677), .B1(N4012), .B2(n2755), .Z(n12196) );
  aor22d1 U1151 ( .A1(n510), .A2(n3677), .B1(N4013), .B2(n2755), .Z(n12197) );
  aor222d1 U1152 ( .A1(N4664), .A2(n3658), .B1(N3915), .B2(n2766), .C1(N4724), 
        .C2(n2), .Z(n12198) );
  oai31d1 U1157 ( .B1(n3667), .B2(new_reference_is_done), .B3(n2775), .A(n3683), .ZN(n12199) );
  aon211d1 U1158 ( .C1(n3670), .C2(n2782), .B(n3667), .A(reading_compare), 
        .ZN(n3683) );
  aon211d1 U1163 ( .C1(n2759), .C2(n3655), .B(n2776), .A(n3686), .ZN(n12200)
         );
  aor22d1 U1166 ( .A1(n513), .A2(n3677), .B1(N5070), .B2(n2755), .Z(n12201) );
  aon211d1 U1168 ( .C1(n3688), .C2(N5285), .B(n3649), .A(n493), .ZN(n3687) );
  oai22d1 U1172 ( .A1(N26480), .A2(n3654), .B1(n3685), .B2(n2774), .ZN(n3689)
         );
  oai21d1 U1175 ( .B1(N5285), .B2(n3676), .A(n2771), .ZN(n3655) );
  oai21d1 U1178 ( .B1(n3690), .B2(n3691), .A(n2772), .ZN(n12203) );
  xr02d1 U1181 ( .A1(count_image[0]), .A2(n963), .Z(n3698) );
  xr02d1 U1182 ( .A1(count_image[1]), .A2(n1034), .Z(n3697) );
  xr02d1 U1183 ( .A1(n2739), .A2(N6870), .Z(n3695) );
  xr02d1 U1184 ( .A1(n2784), .A2(N6869), .Z(n3694) );
  xn02d1 U1185 ( .A1(count_image[6]), .A2(N6873), .ZN(n3693) );
  xr02d1 U1188 ( .A1(\lt_82/A[4] ), .A2(N6871), .Z(n3705) );
  xr02d1 U1189 ( .A1(\lt_82/A[5] ), .A2(N6872), .Z(n3704) );
  xn02d1 U1190 ( .A1(count_image[8]), .A2(N6875), .ZN(n3702) );
  xn02d1 U1192 ( .A1(count_image[7]), .A2(N6874), .ZN(n3701) );
  oai22d1 U1193 ( .A1(n12184), .A2(n497), .B1(n12204), .B2(n3706), .ZN(n12725)
         );
  oai22d1 U1194 ( .A1(n12183), .A2(n497), .B1(n12205), .B2(n3706), .ZN(n12726)
         );
  oai22d1 U1195 ( .A1(n12182), .A2(n497), .B1(n12206), .B2(n3706), .ZN(n12727)
         );
  oai22d1 U1196 ( .A1(n12181), .A2(n497), .B1(n12207), .B2(n3706), .ZN(n12728)
         );
  oai22d1 U1197 ( .A1(n12180), .A2(n497), .B1(n12208), .B2(n3706), .ZN(n12729)
         );
  oai22d1 U1198 ( .A1(n12179), .A2(n497), .B1(n12209), .B2(n3706), .ZN(n12730)
         );
  oai22d1 U1199 ( .A1(n12178), .A2(n497), .B1(n12210), .B2(n3706), .ZN(n12731)
         );
  oai22d1 U1200 ( .A1(n12177), .A2(n497), .B1(n12211), .B2(n3706), .ZN(n12732)
         );
  oai22d1 U1201 ( .A1(n12174), .A2(n497), .B1(n12212), .B2(n3706), .ZN(n12733)
         );
  aor22d1 U1206 ( .A1(N6844), .A2(n3707), .B1(count_image[7]), .B2(n2758), .Z(
        n12734) );
  aor22d1 U1207 ( .A1(N6843), .A2(n3707), .B1(count_image[6]), .B2(n2758), .Z(
        n12735) );
  oaim22d1 U1208 ( .A1(n3707), .A2(n12187), .B1(N6842), .B2(n3707), .ZN(n12736) );
  oaim22d1 U1209 ( .A1(n3707), .A2(n12188), .B1(N6841), .B2(n3707), .ZN(n12737) );
  oaim22d1 U1210 ( .A1(n2739), .A2(n3707), .B1(N6840), .B2(n3707), .ZN(n12738)
         );
  oaim22d1 U1211 ( .A1(n2784), .A2(n3707), .B1(N6839), .B2(n3707), .ZN(n12739)
         );
  aor22d1 U1212 ( .A1(N6838), .A2(n3707), .B1(count_image[1]), .B2(n2758), .Z(
        n12740) );
  aor22d1 U1213 ( .A1(N6837), .A2(n3707), .B1(count_image[0]), .B2(n2758), .Z(
        n12741) );
  aor22d1 U1214 ( .A1(N6845), .A2(n3707), .B1(count_image[8]), .B2(n2758), .Z(
        n12742) );
  oai21d1 U1215 ( .B1(n3709), .B2(n945), .A(n12162), .ZN(n12743) );
  oai21d1 U1216 ( .B1(n945), .B2(n3711), .A(n2809), .ZN(n12744) );
  oai21d1 U1217 ( .B1(n945), .B2(n3713), .A(n12152), .ZN(n12745) );
  oai21d1 U1218 ( .B1(n945), .B2(n3714), .A(n4886), .ZN(n12746) );
  oai21d1 U1219 ( .B1(n945), .B2(n3716), .A(n6654), .ZN(n12747) );
  oai21d1 U1220 ( .B1(n945), .B2(n3718), .A(n5320), .ZN(n12748) );
  oai21d1 U1221 ( .B1(n945), .B2(n3720), .A(n6979), .ZN(n12749) );
  oai21d1 U1222 ( .B1(n945), .B2(n3722), .A(n5797), .ZN(n12750) );
  oai21d1 U1223 ( .B1(n945), .B2(n3724), .A(n6209), .ZN(n12751) );
  oai21d1 U1224 ( .B1(n946), .B2(n3726), .A(n12173), .ZN(n12752) );
  oai21d1 U1225 ( .B1(n946), .B2(n3727), .A(n6508), .ZN(n12753) );
  oai21d1 U1226 ( .B1(n946), .B2(n3729), .A(n4980), .ZN(n12754) );
  oai21d1 U1227 ( .B1(n946), .B2(n3731), .A(n6723), .ZN(n12755) );
  oai21d1 U1228 ( .B1(n946), .B2(n3733), .A(n5470), .ZN(n12756) );
  oai21d1 U1229 ( .B1(n946), .B2(n3735), .A(n7050), .ZN(n12757) );
  oai21d1 U1230 ( .B1(n946), .B2(n3737), .A(n5894), .ZN(n12758) );
  oai21d1 U1231 ( .B1(n946), .B2(n3739), .A(n6276), .ZN(n12759) );
  oai21d1 U1232 ( .B1(n946), .B2(n3741), .A(n4393), .ZN(n12760) );
  oai21d1 U1233 ( .B1(n947), .B2(n3743), .A(n6553), .ZN(n12761) );
  oai21d1 U1234 ( .B1(n947), .B2(n3745), .A(n5118), .ZN(n12762) );
  oai21d1 U1235 ( .B1(n947), .B2(n3747), .A(n6817), .ZN(n12763) );
  oai21d1 U1236 ( .B1(n947), .B2(n3749), .A(n12166), .ZN(n12764) );
  oai21d1 U1237 ( .B1(n947), .B2(n3750), .A(n7115), .ZN(n12765) );
  oai21d1 U1238 ( .B1(n947), .B2(n3752), .A(n5968), .ZN(n12766) );
  oai21d1 U1239 ( .B1(n947), .B2(n3754), .A(n6356), .ZN(n12767) );
  oai21d1 U1240 ( .B1(n947), .B2(n3756), .A(n4633), .ZN(n12768) );
  oai21d1 U1241 ( .B1(n947), .B2(n3758), .A(n6596), .ZN(n12769) );
  oai21d1 U1243 ( .B1(n948), .B2(n3760), .A(n5221), .ZN(n12770) );
  oai21d1 U1244 ( .B1(n948), .B2(n3762), .A(n12125), .ZN(n12771) );
  oai21d1 U1245 ( .B1(n948), .B2(n3763), .A(n5715), .ZN(n12772) );
  oai21d1 U1246 ( .B1(n948), .B2(n3765), .A(n7188), .ZN(n12773) );
  oai21d1 U1247 ( .B1(n944), .B2(n3768), .A(n6074), .ZN(n12774) );
  oai21d1 U1248 ( .B1(n3709), .B2(n944), .A(n12161), .ZN(n12775) );
  oai21d1 U1249 ( .B1(n3711), .B2(n944), .A(n2819), .ZN(n12776) );
  oai21d1 U1250 ( .B1(n3713), .B2(n944), .A(n12151), .ZN(n12777) );
  oai21d1 U1251 ( .B1(n3714), .B2(n944), .A(n4890), .ZN(n12778) );
  oai21d1 U1252 ( .B1(n3716), .B2(n943), .A(n6655), .ZN(n12779) );
  oai21d1 U1253 ( .B1(n3718), .B2(n943), .A(n5322), .ZN(n12780) );
  oai21d1 U1254 ( .B1(n3720), .B2(n943), .A(n6982), .ZN(n12781) );
  oai21d1 U1255 ( .B1(n3722), .B2(n943), .A(n5798), .ZN(n12782) );
  oai21d1 U1256 ( .B1(n3724), .B2(n943), .A(n12158), .ZN(n12783) );
  oai21d1 U1257 ( .B1(n3726), .B2(n943), .A(n4298), .ZN(n12784) );
  oai21d1 U1258 ( .B1(n3727), .B2(n943), .A(n12147), .ZN(n12785) );
  oai21d1 U1259 ( .B1(n3729), .B2(n943), .A(n4984), .ZN(n12786) );
  oai21d1 U1260 ( .B1(n3731), .B2(n943), .A(n6731), .ZN(n12787) );
  oai21d1 U1261 ( .B1(n3733), .B2(n942), .A(n5484), .ZN(n12788) );
  oai21d1 U1262 ( .B1(n3735), .B2(n942), .A(n7057), .ZN(n12789) );
  oai21d1 U1263 ( .B1(n3737), .B2(n942), .A(n5898), .ZN(n12790) );
  oai21d1 U1265 ( .B1(n3739), .B2(n942), .A(n12156), .ZN(n12791) );
  oai21d1 U1266 ( .B1(n3741), .B2(n942), .A(n4397), .ZN(n12792) );
  oai21d1 U1267 ( .B1(n3743), .B2(n942), .A(n6555), .ZN(n12793) );
  oai21d1 U1268 ( .B1(n3745), .B2(n942), .A(n5126), .ZN(n12794) );
  oai21d1 U1269 ( .B1(n3747), .B2(n942), .A(n12129), .ZN(n12795) );
  oai21d1 U1270 ( .B1(n3749), .B2(n942), .A(n5607), .ZN(n12796) );
  oai21d1 U1271 ( .B1(n3750), .B2(n941), .A(n7117), .ZN(n12797) );
  oai21d1 U1272 ( .B1(n3752), .B2(n941), .A(n5979), .ZN(n12798) );
  oai21d1 U1273 ( .B1(n3754), .B2(n941), .A(n6358), .ZN(n12799) );
  oai21d1 U1274 ( .B1(n3756), .B2(n941), .A(n4635), .ZN(n12800) );
  oai21d1 U1275 ( .B1(n3758), .B2(n941), .A(n12141), .ZN(n12801) );
  oai21d1 U1276 ( .B1(n3760), .B2(n941), .A(n5231), .ZN(n12802) );
  oai21d1 U1277 ( .B1(n3762), .B2(n941), .A(n6894), .ZN(n12803) );
  oai21d1 U1278 ( .B1(n3763), .B2(n941), .A(n5727), .ZN(n12804) );
  oai21d1 U1279 ( .B1(n3765), .B2(n941), .A(n7194), .ZN(n12805) );
  oai21d1 U1281 ( .B1(n3768), .B2(n940), .A(n6083), .ZN(n12806) );
  oai21d1 U1282 ( .B1(n3709), .B2(n940), .A(n12160), .ZN(n12807) );
  oai21d1 U1283 ( .B1(n3711), .B2(n940), .A(n2915), .ZN(n12808) );
  oai21d1 U1284 ( .B1(n3713), .B2(n940), .A(n6428), .ZN(n12809) );
  oai21d1 U1285 ( .B1(n3714), .B2(n940), .A(n4894), .ZN(n12810) );
  oai21d1 U1286 ( .B1(n3716), .B2(n939), .A(n6658), .ZN(n12811) );
  oai21d1 U1287 ( .B1(n3718), .B2(n939), .A(n12167), .ZN(n12812) );
  oai21d1 U1288 ( .B1(n3720), .B2(n939), .A(n6990), .ZN(n12813) );
  oai21d1 U1289 ( .B1(n3722), .B2(n939), .A(n5802), .ZN(n12814) );
  oai21d1 U1290 ( .B1(n3724), .B2(n939), .A(n6218), .ZN(n12815) );
  oai21d1 U1291 ( .B1(n3726), .B2(n939), .A(n4300), .ZN(n12816) );
  oai21d1 U1292 ( .B1(n3727), .B2(n939), .A(n6519), .ZN(n12817) );
  oai21d1 U1293 ( .B1(n3729), .B2(n939), .A(n5003), .ZN(n12818) );
  oai21d1 U1294 ( .B1(n3731), .B2(n939), .A(n6732), .ZN(n12819) );
  oai21d1 U1296 ( .B1(n3733), .B2(n938), .A(n5494), .ZN(n12820) );
  oai21d1 U1297 ( .B1(n3735), .B2(n938), .A(n12119), .ZN(n12821) );
  oai21d1 U1298 ( .B1(n3737), .B2(n938), .A(n5902), .ZN(n12822) );
  oai21d1 U1299 ( .B1(n3739), .B2(n938), .A(n6287), .ZN(n12823) );
  oai21d1 U1300 ( .B1(n3741), .B2(n938), .A(n4406), .ZN(n12824) );
  oai21d1 U1301 ( .B1(n3743), .B2(n938), .A(n12142), .ZN(n12825) );
  oai21d1 U1302 ( .B1(n3745), .B2(n938), .A(n5136), .ZN(n12826) );
  oai21d1 U1303 ( .B1(n3747), .B2(n938), .A(n6826), .ZN(n12827) );
  oai21d1 U1304 ( .B1(n3749), .B2(n938), .A(n5617), .ZN(n12828) );
  oai21d1 U1305 ( .B1(n3750), .B2(n937), .A(n7121), .ZN(n12829) );
  oai21d1 U1306 ( .B1(n3752), .B2(n937), .A(n5980), .ZN(n12830) );
  oai21d1 U1307 ( .B1(n3754), .B2(n937), .A(n6360), .ZN(n12831) );
  oai21d1 U1308 ( .B1(n3756), .B2(n937), .A(n4640), .ZN(n12832) );
  oai21d1 U1309 ( .B1(n3758), .B2(n937), .A(n12140), .ZN(n12833) );
  oai21d1 U1310 ( .B1(n3760), .B2(n937), .A(n5235), .ZN(n12834) );
  oai21d1 U1311 ( .B1(n3762), .B2(n937), .A(n6897), .ZN(n12835) );
  oai21d1 U1313 ( .B1(n3763), .B2(n937), .A(n5728), .ZN(n12836) );
  oai21d1 U1314 ( .B1(n3765), .B2(n937), .A(n7205), .ZN(n12837) );
  oai21d1 U1316 ( .B1(n3768), .B2(n936), .A(n6084), .ZN(n12838) );
  oai21d1 U1317 ( .B1(n3709), .B2(n936), .A(n6160), .ZN(n12839) );
  oai21d1 U1318 ( .B1(n3711), .B2(n936), .A(n3129), .ZN(n12840) );
  oai21d1 U1319 ( .B1(n3713), .B2(n936), .A(n12150), .ZN(n12841) );
  oai21d1 U1320 ( .B1(n3714), .B2(n936), .A(n4900), .ZN(n12842) );
  oai21d1 U1321 ( .B1(n3716), .B2(n935), .A(n12136), .ZN(n12843) );
  oai21d1 U1322 ( .B1(n3718), .B2(n935), .A(n5355), .ZN(n12844) );
  oai21d1 U1323 ( .B1(n3720), .B2(n935), .A(n6993), .ZN(n12845) );
  oai21d1 U1324 ( .B1(n3722), .B2(n935), .A(n5806), .ZN(n12846) );
  oai21d1 U1325 ( .B1(n3724), .B2(n935), .A(n6225), .ZN(n12847) );
  oai21d1 U1326 ( .B1(n3726), .B2(n935), .A(n4302), .ZN(n12848) );
  oai21d1 U1327 ( .B1(n3727), .B2(n935), .A(n6523), .ZN(n12849) );
  oai21d1 U1329 ( .B1(n3729), .B2(n935), .A(n5034), .ZN(n12850) );
  oai21d1 U1330 ( .B1(n3731), .B2(n935), .A(n6736), .ZN(n12851) );
  oai21d1 U1331 ( .B1(n3733), .B2(n934), .A(n5506), .ZN(n12852) );
  oai21d1 U1332 ( .B1(n3735), .B2(n934), .A(n7066), .ZN(n12853) );
  oai21d1 U1333 ( .B1(n3737), .B2(n934), .A(n5906), .ZN(n12854) );
  oai21d1 U1334 ( .B1(n3739), .B2(n934), .A(n6291), .ZN(n12855) );
  oai21d1 U1335 ( .B1(n3741), .B2(n934), .A(n12171), .ZN(n12856) );
  oai21d1 U1336 ( .B1(n3743), .B2(n934), .A(n6558), .ZN(n12857) );
  oai21d1 U1337 ( .B1(n3745), .B2(n934), .A(n5145), .ZN(n12858) );
  oai21d1 U1338 ( .B1(n3747), .B2(n934), .A(n6837), .ZN(n12859) );
  oai21d1 U1339 ( .B1(n3749), .B2(n934), .A(n5625), .ZN(n12860) );
  oai21d1 U1340 ( .B1(n3750), .B2(n933), .A(n7127), .ZN(n12861) );
  oai21d1 U1341 ( .B1(n3752), .B2(n933), .A(n5982), .ZN(n12862) );
  oai21d1 U1342 ( .B1(n3754), .B2(n933), .A(n6366), .ZN(n12863) );
  oai21d1 U1343 ( .B1(n3756), .B2(n933), .A(n4649), .ZN(n12864) );
  oai21d1 U1344 ( .B1(n3758), .B2(n933), .A(n12139), .ZN(n12865) );
  oai21d1 U1345 ( .B1(n3760), .B2(n933), .A(n5242), .ZN(n12866) );
  oai21d1 U1346 ( .B1(n3762), .B2(n933), .A(n12124), .ZN(n12867) );
  oai21d1 U1347 ( .B1(n3763), .B2(n933), .A(n5730), .ZN(n12868) );
  oai21d1 U1348 ( .B1(n3765), .B2(n933), .A(n7207), .ZN(n12869) );
  oai21d1 U1351 ( .B1(n3768), .B2(n932), .A(n6089), .ZN(n12870) );
  oai21d1 U1352 ( .B1(n3709), .B2(n932), .A(n6162), .ZN(n12871) );
  oai21d1 U1353 ( .B1(n3711), .B2(n932), .A(n3138), .ZN(n12872) );
  oai21d1 U1354 ( .B1(n3713), .B2(n932), .A(n6443), .ZN(n12873) );
  oai21d1 U1356 ( .B1(n3714), .B2(n932), .A(n4902), .ZN(n12874) );
  oai21d1 U1357 ( .B1(n3716), .B2(n931), .A(n12135), .ZN(n12875) );
  oai21d1 U1358 ( .B1(n3718), .B2(n931), .A(n5370), .ZN(n12876) );
  oai21d1 U1359 ( .B1(n3720), .B2(n931), .A(n6997), .ZN(n12877) );
  oai21d1 U1360 ( .B1(n3722), .B2(n931), .A(n5818), .ZN(n12878) );
  oai21d1 U1361 ( .B1(n3724), .B2(n931), .A(n6229), .ZN(n12879) );
  oai21d1 U1362 ( .B1(n3726), .B2(n931), .A(n4304), .ZN(n12880) );
  oai21d1 U1363 ( .B1(n3727), .B2(n931), .A(n6525), .ZN(n12881) );
  oai21d1 U1364 ( .B1(n3729), .B2(n931), .A(n5043), .ZN(n12882) );
  oai21d1 U1365 ( .B1(n3731), .B2(n931), .A(n12132), .ZN(n12883) );
  oai21d1 U1366 ( .B1(n3733), .B2(n930), .A(n5523), .ZN(n12884) );
  oai21d1 U1367 ( .B1(n3735), .B2(n930), .A(n7067), .ZN(n12885) );
  oai21d1 U1368 ( .B1(n3737), .B2(n930), .A(n5920), .ZN(n12886) );
  oai21d1 U1369 ( .B1(n3739), .B2(n930), .A(n6293), .ZN(n12887) );
  oai21d1 U1370 ( .B1(n3741), .B2(n930), .A(n4419), .ZN(n12888) );
  oai21d1 U1371 ( .B1(n3743), .B2(n930), .A(n6560), .ZN(n12889) );
  oai21d1 U1373 ( .B1(n3745), .B2(n930), .A(n5146), .ZN(n12890) );
  oai21d1 U1374 ( .B1(n3747), .B2(n930), .A(n6838), .ZN(n12891) );
  oai21d1 U1375 ( .B1(n3749), .B2(n930), .A(n12165), .ZN(n12892) );
  oai21d1 U1376 ( .B1(n3750), .B2(n929), .A(n7133), .ZN(n12893) );
  oai21d1 U1377 ( .B1(n3752), .B2(n929), .A(n5988), .ZN(n12894) );
  oai21d1 U1378 ( .B1(n3754), .B2(n929), .A(n6368), .ZN(n12895) );
  oai21d1 U1379 ( .B1(n3756), .B2(n929), .A(n4653), .ZN(n12896) );
  oai21d1 U1380 ( .B1(n3758), .B2(n929), .A(n12138), .ZN(n12897) );
  oai21d1 U1381 ( .B1(n3760), .B2(n929), .A(n5249), .ZN(n12898) );
  oai21d1 U1382 ( .B1(n3762), .B2(n929), .A(n12123), .ZN(n12899) );
  oai21d1 U1383 ( .B1(n3763), .B2(n929), .A(n5732), .ZN(n12900) );
  oai21d1 U1384 ( .B1(n3765), .B2(n929), .A(n7222), .ZN(n12901) );
  oai21d1 U1386 ( .B1(n3768), .B2(n928), .A(n6097), .ZN(n12902) );
  oai21d1 U1387 ( .B1(n3709), .B2(n928), .A(n6166), .ZN(n12903) );
  oai21d1 U1388 ( .B1(n3711), .B2(n928), .A(n3268), .ZN(n12904) );
  oai21d1 U1389 ( .B1(n3713), .B2(n928), .A(n6445), .ZN(n12905) );
  oai21d1 U1390 ( .B1(n3714), .B2(n928), .A(n4915), .ZN(n12906) );
  oai21d1 U1391 ( .B1(n3716), .B2(n927), .A(n6670), .ZN(n12907) );
  oai21d1 U1392 ( .B1(n3718), .B2(n927), .A(n5397), .ZN(n12908) );
  oai21d1 U1393 ( .B1(n3720), .B2(n927), .A(n6998), .ZN(n12909) );
  oai21d1 U1394 ( .B1(n3722), .B2(n927), .A(n5825), .ZN(n12910) );
  oai21d1 U1395 ( .B1(n3724), .B2(n927), .A(n12157), .ZN(n12911) );
  oai21d1 U1396 ( .B1(n3726), .B2(n927), .A(n4306), .ZN(n12912) );
  oai21d1 U1397 ( .B1(n3727), .B2(n927), .A(n6529), .ZN(n12913) );
  oai21d1 U1398 ( .B1(n3729), .B2(n927), .A(n5046), .ZN(n12914) );
  oai21d1 U1399 ( .B1(n3731), .B2(n927), .A(n6747), .ZN(n12915) );
  oai21d1 U1400 ( .B1(n3733), .B2(n926), .A(n5527), .ZN(n12916) );
  oai21d1 U1401 ( .B1(n3735), .B2(n926), .A(n7069), .ZN(n12917) );
  oai21d1 U1402 ( .B1(n3737), .B2(n926), .A(n5927), .ZN(n12918) );
  oai21d1 U1403 ( .B1(n3739), .B2(n926), .A(n6297), .ZN(n12919) );
  oai21d1 U1404 ( .B1(n3741), .B2(n926), .A(n4427), .ZN(n12920) );
  oai21d1 U1405 ( .B1(n3743), .B2(n926), .A(n6562), .ZN(n12921) );
  oai21d1 U1406 ( .B1(n3745), .B2(n926), .A(n5156), .ZN(n12922) );
  oai21d1 U1407 ( .B1(n3747), .B2(n926), .A(n6840), .ZN(n12923) );
  oai21d1 U1408 ( .B1(n3749), .B2(n926), .A(n5633), .ZN(n12924) );
  oai21d1 U1409 ( .B1(n3750), .B2(n925), .A(n7136), .ZN(n12925) );
  oai21d1 U1410 ( .B1(n3752), .B2(n925), .A(n6004), .ZN(n12926) );
  oai21d1 U1411 ( .B1(n3754), .B2(n925), .A(n6371), .ZN(n12927) );
  oai21d1 U1412 ( .B1(n3756), .B2(n925), .A(n4663), .ZN(n12928) );
  oai21d1 U1413 ( .B1(n3758), .B2(n925), .A(n6606), .ZN(n12929) );
  oai21d1 U1414 ( .B1(n3760), .B2(n925), .A(n5254), .ZN(n12930) );
  oai21d1 U1415 ( .B1(n3762), .B2(n925), .A(n6919), .ZN(n12931) );
  oai21d1 U1416 ( .B1(n3763), .B2(n925), .A(n5737), .ZN(n12932) );
  oai21d1 U1417 ( .B1(n3765), .B2(n925), .A(n7232), .ZN(n12933) );
  oai21d1 U1419 ( .B1(n3768), .B2(n924), .A(n6098), .ZN(n12934) );
  oai21d1 U1420 ( .B1(n3709), .B2(n924), .A(n6170), .ZN(n12935) );
  oai21d1 U1421 ( .B1(n3711), .B2(n924), .A(n3331), .ZN(n12936) );
  oai21d1 U1422 ( .B1(n3713), .B2(n924), .A(n6455), .ZN(n12937) );
  oai21d1 U1423 ( .B1(n3714), .B2(n924), .A(n4939), .ZN(n12938) );
  oai21d1 U1424 ( .B1(n3716), .B2(n923), .A(n6675), .ZN(n12939) );
  oai21d1 U1425 ( .B1(n3718), .B2(n923), .A(n5405), .ZN(n12940) );
  oai21d1 U1426 ( .B1(n3720), .B2(n923), .A(n7006), .ZN(n12941) );
  oai21d1 U1427 ( .B1(n3722), .B2(n923), .A(n5826), .ZN(n12942) );
  oai21d1 U1428 ( .B1(n3724), .B2(n923), .A(n6240), .ZN(n12943) );
  oai21d1 U1429 ( .B1(n3726), .B2(n923), .A(n4307), .ZN(n12944) );
  oai21d1 U1430 ( .B1(n3727), .B2(n923), .A(n12146), .ZN(n12945) );
  oai21d1 U1431 ( .B1(n3729), .B2(n923), .A(n5049), .ZN(n12946) );
  oai21d1 U1432 ( .B1(n3731), .B2(n923), .A(n6752), .ZN(n12947) );
  oai21d1 U1433 ( .B1(n3733), .B2(n922), .A(n5531), .ZN(n12948) );
  oai21d1 U1434 ( .B1(n3735), .B2(n922), .A(n7072), .ZN(n12949) );
  oai21d1 U1435 ( .B1(n3737), .B2(n922), .A(n5931), .ZN(n12950) );
  oai21d1 U1436 ( .B1(n3739), .B2(n922), .A(n6303), .ZN(n12951) );
  oai21d1 U1437 ( .B1(n3741), .B2(n922), .A(n4436), .ZN(n12952) );
  oai21d1 U1438 ( .B1(n3743), .B2(n922), .A(n6565), .ZN(n12953) );
  oai21d1 U1439 ( .B1(n3745), .B2(n922), .A(n5164), .ZN(n12954) );
  oai21d1 U1440 ( .B1(n3747), .B2(n922), .A(n6842), .ZN(n12955) );
  oai21d1 U1441 ( .B1(n3749), .B2(n922), .A(n5636), .ZN(n12956) );
  oai21d1 U1442 ( .B1(n3750), .B2(n921), .A(n7150), .ZN(n12957) );
  oai21d1 U1443 ( .B1(n3752), .B2(n921), .A(n6007), .ZN(n12958) );
  oai21d1 U1444 ( .B1(n3754), .B2(n921), .A(n12153), .ZN(n12959) );
  oai21d1 U1445 ( .B1(n3756), .B2(n921), .A(n4675), .ZN(n12960) );
  oai21d1 U1446 ( .B1(n3758), .B2(n921), .A(n6613), .ZN(n12961) );
  oai21d1 U1447 ( .B1(n3760), .B2(n921), .A(n5265), .ZN(n12962) );
  oai21d1 U1448 ( .B1(n3762), .B2(n921), .A(n12122), .ZN(n12963) );
  oai21d1 U1449 ( .B1(n3763), .B2(n921), .A(n5738), .ZN(n12964) );
  oai21d1 U1450 ( .B1(n3765), .B2(n921), .A(n7237), .ZN(n12965) );
  oai21d1 U1452 ( .B1(n3768), .B2(n920), .A(n6100), .ZN(n12966) );
  oai21d1 U1453 ( .B1(n3709), .B2(n920), .A(n6173), .ZN(n12967) );
  oai21d1 U1454 ( .B1(n3711), .B2(n920), .A(n3478), .ZN(n12968) );
  oai21d1 U1455 ( .B1(n3713), .B2(n920), .A(n12149), .ZN(n12969) );
  oai21d1 U1456 ( .B1(n3714), .B2(n920), .A(n12169), .ZN(n12970) );
  oai21d1 U1457 ( .B1(n3716), .B2(n919), .A(n6676), .ZN(n12971) );
  oai21d1 U1459 ( .B1(n3718), .B2(n919), .A(n5410), .ZN(n12972) );
  oai21d1 U1460 ( .B1(n3720), .B2(n919), .A(n7016), .ZN(n12973) );
  oai21d1 U1461 ( .B1(n3722), .B2(n919), .A(n5834), .ZN(n12974) );
  oai21d1 U1462 ( .B1(n3724), .B2(n919), .A(n6242), .ZN(n12975) );
  oai21d1 U1463 ( .B1(n3726), .B2(n919), .A(n4311), .ZN(n12976) );
  oai21d1 U1464 ( .B1(n3727), .B2(n919), .A(n6533), .ZN(n12977) );
  oai21d1 U1465 ( .B1(n3729), .B2(n919), .A(n5060), .ZN(n12978) );
  oai21d1 U1466 ( .B1(n3731), .B2(n919), .A(n6753), .ZN(n12979) );
  oai21d1 U1467 ( .B1(n3733), .B2(n918), .A(n5540), .ZN(n12980) );
  oai21d1 U1468 ( .B1(n3735), .B2(n918), .A(n7075), .ZN(n12981) );
  oai21d1 U1469 ( .B1(n3737), .B2(n918), .A(n5933), .ZN(n12982) );
  oai21d1 U1470 ( .B1(n3739), .B2(n918), .A(n6305), .ZN(n12983) );
  oai21d1 U1471 ( .B1(n3741), .B2(n918), .A(n4450), .ZN(n12984) );
  oai21d1 U1472 ( .B1(n3743), .B2(n918), .A(n6566), .ZN(n12985) );
  oai21d1 U1473 ( .B1(n3745), .B2(n918), .A(n5168), .ZN(n12986) );
  oai21d1 U1474 ( .B1(n3747), .B2(n918), .A(n6849), .ZN(n12987) );
  oai21d1 U1475 ( .B1(n3749), .B2(n918), .A(n5644), .ZN(n12988) );
  oai21d1 U1476 ( .B1(n3750), .B2(n917), .A(n7152), .ZN(n12989) );
  oai21d1 U1477 ( .B1(n3752), .B2(n917), .A(n6024), .ZN(n12990) );
  oai21d1 U1478 ( .B1(n3754), .B2(n917), .A(n6388), .ZN(n12991) );
  oai21d1 U1479 ( .B1(n3756), .B2(n917), .A(n4689), .ZN(n12992) );
  oai21d1 U1480 ( .B1(n3758), .B2(n917), .A(n6618), .ZN(n12993) );
  oai21d1 U1481 ( .B1(n3760), .B2(n917), .A(n5266), .ZN(n12994) );
  oai21d1 U1482 ( .B1(n3762), .B2(n917), .A(n6923), .ZN(n12995) );
  oai21d1 U1483 ( .B1(n3763), .B2(n917), .A(n5746), .ZN(n12996) );
  oai21d1 U1484 ( .B1(n3765), .B2(n917), .A(n7240), .ZN(n12997) );
  oai21d1 U1486 ( .B1(n3768), .B2(n916), .A(n6113), .ZN(n12998) );
  oai21d1 U1487 ( .B1(n3709), .B2(n916), .A(n6174), .ZN(n12999) );
  oai21d1 U1488 ( .B1(n3711), .B2(n916), .A(n3577), .ZN(n13000) );
  oai21d1 U1489 ( .B1(n3713), .B2(n916), .A(n6469), .ZN(n13001) );
  oai21d1 U1490 ( .B1(n3714), .B2(n916), .A(n4948), .ZN(n13002) );
  oai21d1 U1491 ( .B1(n3716), .B2(n915), .A(n6677), .ZN(n13003) );
  oai21d1 U1492 ( .B1(n3718), .B2(n915), .A(n5426), .ZN(n13004) );
  oai21d1 U1493 ( .B1(n3720), .B2(n915), .A(n7017), .ZN(n13005) );
  oai21d1 U1494 ( .B1(n3722), .B2(n915), .A(n5835), .ZN(n13006) );
  oai21d1 U1495 ( .B1(n3724), .B2(n915), .A(n6246), .ZN(n13007) );
  oai21d1 U1496 ( .B1(n3726), .B2(n915), .A(n4313), .ZN(n13008) );
  oai21d1 U1497 ( .B1(n3727), .B2(n915), .A(n6538), .ZN(n13009) );
  oai21d1 U1498 ( .B1(n3729), .B2(n915), .A(n5063), .ZN(n13010) );
  oai21d1 U1499 ( .B1(n3731), .B2(n915), .A(n6759), .ZN(n13011) );
  oai21d1 U1500 ( .B1(n3733), .B2(n914), .A(n5542), .ZN(n13012) );
  oai21d1 U1501 ( .B1(n3735), .B2(n914), .A(n7076), .ZN(n13013) );
  oai21d1 U1502 ( .B1(n3737), .B2(n914), .A(n5937), .ZN(n13014) );
  oai21d1 U1503 ( .B1(n3739), .B2(n914), .A(n6310), .ZN(n13015) );
  oai21d1 U1504 ( .B1(n3741), .B2(n914), .A(n4451), .ZN(n13016) );
  oai21d1 U1505 ( .B1(n3743), .B2(n914), .A(n6567), .ZN(n13017) );
  oai21d1 U1506 ( .B1(n3745), .B2(n914), .A(n5173), .ZN(n13018) );
  oai21d1 U1507 ( .B1(n3747), .B2(n914), .A(n6855), .ZN(n13019) );
  oai21d1 U1508 ( .B1(n3749), .B2(n914), .A(n5648), .ZN(n13020) );
  oai21d1 U1509 ( .B1(n3750), .B2(n913), .A(n12118), .ZN(n13021) );
  oai21d1 U1510 ( .B1(n3752), .B2(n913), .A(n6025), .ZN(n13022) );
  oai21d1 U1511 ( .B1(n3754), .B2(n913), .A(n6389), .ZN(n13023) );
  oai21d1 U1512 ( .B1(n3756), .B2(n913), .A(n4691), .ZN(n13024) );
  oai21d1 U1513 ( .B1(n3758), .B2(n913), .A(n12137), .ZN(n13025) );
  oai21d1 U1514 ( .B1(n3760), .B2(n913), .A(n5268), .ZN(n13026) );
  oai21d1 U1515 ( .B1(n3762), .B2(n913), .A(n12121), .ZN(n13027) );
  oai21d1 U1516 ( .B1(n3763), .B2(n913), .A(n5747), .ZN(n13028) );
  oai21d1 U1517 ( .B1(n3765), .B2(n913), .A(n7242), .ZN(n13029) );
  oai21d1 U1519 ( .B1(n3768), .B2(n912), .A(n6115), .ZN(n13030) );
  oai21d1 U1520 ( .B1(n3709), .B2(n912), .A(n6176), .ZN(n13031) );
  oai21d1 U1522 ( .B1(n3711), .B2(n912), .A(n3619), .ZN(n13032) );
  oai21d1 U1523 ( .B1(n3713), .B2(n912), .A(n6475), .ZN(n13033) );
  oai21d1 U1524 ( .B1(n3714), .B2(n912), .A(n4951), .ZN(n13034) );
  oai21d1 U1525 ( .B1(n3716), .B2(n911), .A(n12134), .ZN(n13035) );
  oai21d1 U1526 ( .B1(n3718), .B2(n911), .A(n5431), .ZN(n13036) );
  oai21d1 U1527 ( .B1(n3720), .B2(n911), .A(n7019), .ZN(n13037) );
  oai21d1 U1528 ( .B1(n3722), .B2(n911), .A(n5839), .ZN(n13038) );
  oai21d1 U1529 ( .B1(n3724), .B2(n911), .A(n6250), .ZN(n13039) );
  oai21d1 U1530 ( .B1(n3726), .B2(n911), .A(n4314), .ZN(n13040) );
  oai21d1 U1531 ( .B1(n3727), .B2(n911), .A(n6540), .ZN(n13041) );
  oai21d1 U1532 ( .B1(n3729), .B2(n911), .A(n5068), .ZN(n13042) );
  oai21d1 U1533 ( .B1(n3731), .B2(n911), .A(n6776), .ZN(n13043) );
  oai21d1 U1535 ( .B1(n3733), .B2(n910), .A(n5548), .ZN(n13044) );
  oai21d1 U1536 ( .B1(n3735), .B2(n910), .A(n7079), .ZN(n13045) );
  oai21d1 U1537 ( .B1(n3737), .B2(n910), .A(n5944), .ZN(n13046) );
  oai21d1 U1538 ( .B1(n3739), .B2(n910), .A(n12155), .ZN(n13047) );
  oai21d1 U1539 ( .B1(n3741), .B2(n910), .A(n4459), .ZN(n13048) );
  oai21d1 U1540 ( .B1(n3743), .B2(n910), .A(n6571), .ZN(n13049) );
  oai21d1 U1541 ( .B1(n3745), .B2(n910), .A(n5186), .ZN(n13050) );
  oai21d1 U1542 ( .B1(n3747), .B2(n910), .A(n12128), .ZN(n13051) );
  oai21d1 U1543 ( .B1(n3749), .B2(n910), .A(n5669), .ZN(n13052) );
  oai21d1 U1544 ( .B1(n3750), .B2(n909), .A(n7155), .ZN(n13053) );
  oai21d1 U1545 ( .B1(n3752), .B2(n909), .A(n6038), .ZN(n13054) );
  oai21d1 U1546 ( .B1(n3754), .B2(n909), .A(n6390), .ZN(n13055) );
  oai21d1 U1547 ( .B1(n3756), .B2(n909), .A(n12170), .ZN(n13056) );
  oai21d1 U1548 ( .B1(n3758), .B2(n909), .A(n6628), .ZN(n13057) );
  oai21d1 U1549 ( .B1(n3760), .B2(n909), .A(n5276), .ZN(n13058) );
  oai21d1 U1550 ( .B1(n3762), .B2(n909), .A(n6934), .ZN(n13059) );
  oai21d1 U1551 ( .B1(n3763), .B2(n909), .A(n5749), .ZN(n13060) );
  oai21d1 U1552 ( .B1(n3765), .B2(n909), .A(n7243), .ZN(n13061) );
  oai21d1 U1554 ( .B1(n3768), .B2(n908), .A(n6119), .ZN(n13062) );
  oai21d1 U1555 ( .B1(n3709), .B2(n908), .A(n12159), .ZN(n13063) );
  oai21d1 U1556 ( .B1(n3711), .B2(n908), .A(n3814), .ZN(n13064) );
  oai21d1 U1557 ( .B1(n3713), .B2(n908), .A(n6481), .ZN(n13065) );
  oai21d1 U1558 ( .B1(n3714), .B2(n908), .A(n12168), .ZN(n13066) );
  oai21d1 U1559 ( .B1(n3716), .B2(n907), .A(n6683), .ZN(n13067) );
  oai21d1 U1560 ( .B1(n3718), .B2(n907), .A(n5434), .ZN(n13068) );
  oai21d1 U1561 ( .B1(n3720), .B2(n907), .A(n7022), .ZN(n13069) );
  oai21d1 U1562 ( .B1(n3722), .B2(n907), .A(n5846), .ZN(n13070) );
  oai21d1 U1563 ( .B1(n3724), .B2(n907), .A(n6259), .ZN(n13071) );
  oai21d1 U1564 ( .B1(n3726), .B2(n907), .A(n4316), .ZN(n13072) );
  oai21d1 U1565 ( .B1(n3727), .B2(n907), .A(n12145), .ZN(n13073) );
  oai21d1 U1566 ( .B1(n3729), .B2(n907), .A(n5079), .ZN(n13074) );
  oai21d1 U1567 ( .B1(n3731), .B2(n907), .A(n6777), .ZN(n13075) );
  oai21d1 U1568 ( .B1(n3733), .B2(n906), .A(n5558), .ZN(n13076) );
  oai21d1 U1569 ( .B1(n3735), .B2(n906), .A(n7081), .ZN(n13077) );
  oai21d1 U1570 ( .B1(n3737), .B2(n906), .A(n5949), .ZN(n13078) );
  oai21d1 U1571 ( .B1(n3739), .B2(n906), .A(n12154), .ZN(n13079) );
  oai21d1 U1572 ( .B1(n3741), .B2(n906), .A(n4464), .ZN(n13080) );
  oai21d1 U1573 ( .B1(n3743), .B2(n906), .A(n6572), .ZN(n13081) );
  oai21d1 U1574 ( .B1(n3745), .B2(n906), .A(n5189), .ZN(n13082) );
  oai21d1 U1575 ( .B1(n3747), .B2(n906), .A(n6866), .ZN(n13083) );
  oai21d1 U1576 ( .B1(n3749), .B2(n906), .A(n5676), .ZN(n13084) );
  oai21d1 U1577 ( .B1(n3750), .B2(n905), .A(n7166), .ZN(n13085) );
  oai21d1 U1578 ( .B1(n3752), .B2(n905), .A(n6039), .ZN(n13086) );
  oai21d1 U1579 ( .B1(n3754), .B2(n905), .A(n6395), .ZN(n13087) );
  oai21d1 U1580 ( .B1(n3756), .B2(n905), .A(n4703), .ZN(n13088) );
  oai21d1 U1581 ( .B1(n3758), .B2(n905), .A(n6630), .ZN(n13089) );
  oai21d1 U1582 ( .B1(n3760), .B2(n905), .A(n5278), .ZN(n13090) );
  oai21d1 U1583 ( .B1(n3762), .B2(n905), .A(n6938), .ZN(n13091) );
  oai21d1 U1584 ( .B1(n3763), .B2(n905), .A(n5762), .ZN(n13092) );
  oai21d1 U1585 ( .B1(n3765), .B2(n905), .A(n7244), .ZN(n13093) );
  oai21d1 U1587 ( .B1(n3768), .B2(n904), .A(n6123), .ZN(n13094) );
  oai21d1 U1588 ( .B1(n3709), .B2(n904), .A(n6185), .ZN(n13095) );
  oai21d1 U1589 ( .B1(n3711), .B2(n904), .A(n3903), .ZN(n13096) );
  oai21d1 U1590 ( .B1(n3713), .B2(n904), .A(n6484), .ZN(n13097) );
  oai21d1 U1591 ( .B1(n3714), .B2(n904), .A(n4959), .ZN(n13098) );
  oai21d1 U1592 ( .B1(n3716), .B2(n903), .A(n6693), .ZN(n13099) );
  oai21d1 U1593 ( .B1(n3718), .B2(n903), .A(n5440), .ZN(n13100) );
  oai21d1 U1594 ( .B1(n3720), .B2(n903), .A(n7023), .ZN(n13101) );
  oai21d1 U1595 ( .B1(n3722), .B2(n903), .A(n5851), .ZN(n13102) );
  oai21d1 U1596 ( .B1(n3724), .B2(n903), .A(n6264), .ZN(n13103) );
  oai21d1 U1597 ( .B1(n3726), .B2(n903), .A(n4319), .ZN(n13104) );
  oai21d1 U1598 ( .B1(n3727), .B2(n903), .A(n12144), .ZN(n13105) );
  oai21d1 U1599 ( .B1(n3729), .B2(n903), .A(n5098), .ZN(n13106) );
  oai21d1 U1600 ( .B1(n3731), .B2(n903), .A(n6778), .ZN(n13107) );
  oai21d1 U1601 ( .B1(n3733), .B2(n902), .A(n5573), .ZN(n13108) );
  oai21d1 U1602 ( .B1(n3735), .B2(n902), .A(n7093), .ZN(n13109) );
  oai21d1 U1603 ( .B1(n3737), .B2(n902), .A(n5952), .ZN(n13110) );
  oai21d1 U1604 ( .B1(n3739), .B2(n902), .A(n6330), .ZN(n13111) );
  oai21d1 U1605 ( .B1(n3741), .B2(n902), .A(n4491), .ZN(n13112) );
  oai21d1 U1606 ( .B1(n3743), .B2(n902), .A(n6575), .ZN(n13113) );
  oai21d1 U1607 ( .B1(n3745), .B2(n902), .A(n5194), .ZN(n13114) );
  oai21d1 U1608 ( .B1(n3747), .B2(n902), .A(n12127), .ZN(n13115) );
  oai21d1 U1609 ( .B1(n3749), .B2(n902), .A(n5684), .ZN(n13116) );
  oai21d1 U1610 ( .B1(n3750), .B2(n901), .A(n7173), .ZN(n13117) );
  oai21d1 U1611 ( .B1(n3752), .B2(n901), .A(n6051), .ZN(n13118) );
  oai21d1 U1612 ( .B1(n3754), .B2(n901), .A(n6397), .ZN(n13119) );
  oai21d1 U1613 ( .B1(n3756), .B2(n901), .A(n4727), .ZN(n13120) );
  oai21d1 U1615 ( .B1(n3758), .B2(n901), .A(n6638), .ZN(n13121) );
  oai21d1 U1617 ( .B1(n3760), .B2(n901), .A(n5281), .ZN(n13122) );
  oai21d1 U1618 ( .B1(n3762), .B2(n901), .A(n6946), .ZN(n13123) );
  oai21d1 U1619 ( .B1(n3763), .B2(n901), .A(n5768), .ZN(n13124) );
  oai21d1 U1620 ( .B1(n3765), .B2(n901), .A(n7245), .ZN(n13125) );
  oai21d1 U1624 ( .B1(n3768), .B2(n900), .A(n6133), .ZN(n13126) );
  oai21d1 U1625 ( .B1(n3709), .B2(n900), .A(n6189), .ZN(n13127) );
  oai21d1 U1626 ( .B1(n3711), .B2(n900), .A(n3986), .ZN(n13128) );
  oai21d1 U1627 ( .B1(n3713), .B2(n900), .A(n6488), .ZN(n13129) );
  oai21d1 U1628 ( .B1(n3714), .B2(n900), .A(n4965), .ZN(n13130) );
  oai21d1 U1629 ( .B1(n3716), .B2(n899), .A(n6698), .ZN(n13131) );
  oai21d1 U1631 ( .B1(n3718), .B2(n899), .A(n5447), .ZN(n13132) );
  oai21d1 U1632 ( .B1(n3720), .B2(n899), .A(n7034), .ZN(n13133) );
  oai21d1 U1633 ( .B1(n3722), .B2(n899), .A(n5855), .ZN(n13134) );
  oai21d1 U1634 ( .B1(n3724), .B2(n899), .A(n6267), .ZN(n13135) );
  oai21d1 U1635 ( .B1(n3726), .B2(n899), .A(n4321), .ZN(n13136) );
  oai21d1 U1636 ( .B1(n3727), .B2(n899), .A(n12143), .ZN(n13137) );
  oai21d1 U1637 ( .B1(n3729), .B2(n899), .A(n5104), .ZN(n13138) );
  oai21d1 U1638 ( .B1(n3731), .B2(n899), .A(n12131), .ZN(n13139) );
  oai21d1 U1639 ( .B1(n3733), .B2(n898), .A(n5575), .ZN(n13140) );
  oai21d1 U1640 ( .B1(n3735), .B2(n898), .A(n7097), .ZN(n13141) );
  oai21d1 U1641 ( .B1(n3737), .B2(n898), .A(n5957), .ZN(n13142) );
  oai21d1 U1642 ( .B1(n3739), .B2(n898), .A(n6344), .ZN(n13143) );
  oai21d1 U1643 ( .B1(n3741), .B2(n898), .A(n4493), .ZN(n13144) );
  oai21d1 U1644 ( .B1(n3743), .B2(n898), .A(n6576), .ZN(n13145) );
  oai21d1 U1645 ( .B1(n3745), .B2(n898), .A(n5203), .ZN(n13146) );
  oai21d1 U1646 ( .B1(n3747), .B2(n898), .A(n6875), .ZN(n13147) );
  oai21d1 U1647 ( .B1(n3749), .B2(n898), .A(n5689), .ZN(n13148) );
  oai21d1 U1648 ( .B1(n3750), .B2(n897), .A(n7176), .ZN(n13149) );
  oai21d1 U1649 ( .B1(n3752), .B2(n897), .A(n6056), .ZN(n13150) );
  oai21d1 U1650 ( .B1(n3754), .B2(n897), .A(n6400), .ZN(n13151) );
  oai21d1 U1651 ( .B1(n3756), .B2(n897), .A(n4745), .ZN(n13152) );
  oai21d1 U1652 ( .B1(n3758), .B2(n897), .A(n6639), .ZN(n13153) );
  oai21d1 U1653 ( .B1(n3760), .B2(n897), .A(n5284), .ZN(n13154) );
  oai21d1 U1654 ( .B1(n3762), .B2(n897), .A(n6948), .ZN(n13155) );
  oai21d1 U1655 ( .B1(n3763), .B2(n897), .A(n5775), .ZN(n13156) );
  oai21d1 U1656 ( .B1(n3765), .B2(n897), .A(n7251), .ZN(n13157) );
  oai21d1 U1658 ( .B1(n3768), .B2(n896), .A(n6138), .ZN(n13158) );
  oai21d1 U1659 ( .B1(n3709), .B2(n896), .A(n6199), .ZN(n13159) );
  oai21d1 U1661 ( .B1(n3711), .B2(n896), .A(n4119), .ZN(n13160) );
  oai21d1 U1662 ( .B1(n3713), .B2(n896), .A(n12148), .ZN(n13161) );
  oai21d1 U1663 ( .B1(n3714), .B2(n896), .A(n4973), .ZN(n13162) );
  oai21d1 U1664 ( .B1(n3716), .B2(n895), .A(n12133), .ZN(n13163) );
  oai21d1 U1665 ( .B1(n3718), .B2(n895), .A(n5456), .ZN(n13164) );
  oai21d1 U1666 ( .B1(n3720), .B2(n895), .A(n7042), .ZN(n13165) );
  oai21d1 U1667 ( .B1(n3722), .B2(n895), .A(n5858), .ZN(n13166) );
  oai21d1 U1668 ( .B1(n3724), .B2(n895), .A(n6268), .ZN(n13167) );
  oai21d1 U1669 ( .B1(n3726), .B2(n895), .A(n4326), .ZN(n13168) );
  oai21d1 U1670 ( .B1(n3727), .B2(n895), .A(n6548), .ZN(n13169) );
  oai21d1 U1671 ( .B1(n3729), .B2(n895), .A(n5106), .ZN(n13170) );
  oai21d1 U1672 ( .B1(n3731), .B2(n895), .A(n6805), .ZN(n13171) );
  oai21d1 U1673 ( .B1(n3733), .B2(n894), .A(n5581), .ZN(n13172) );
  oai21d1 U1674 ( .B1(n3735), .B2(n894), .A(n7104), .ZN(n13173) );
  oai21d1 U1675 ( .B1(n3737), .B2(n894), .A(n5958), .ZN(n13174) );
  oai21d1 U1676 ( .B1(n3739), .B2(n894), .A(n6345), .ZN(n13175) );
  oai21d1 U1677 ( .B1(n3741), .B2(n894), .A(n4503), .ZN(n13176) );
  oai21d1 U1678 ( .B1(n3743), .B2(n894), .A(n6586), .ZN(n13177) );
  oai21d1 U1679 ( .B1(n3745), .B2(n894), .A(n5204), .ZN(n13178) );
  oai21d1 U1680 ( .B1(n3747), .B2(n894), .A(n6882), .ZN(n13179) );
  oai21d1 U1681 ( .B1(n3749), .B2(n894), .A(n5691), .ZN(n13180) );
  oai21d1 U1682 ( .B1(n3750), .B2(n893), .A(n7182), .ZN(n13181) );
  oai21d1 U1683 ( .B1(n3752), .B2(n893), .A(n6061), .ZN(n13182) );
  oai21d1 U1684 ( .B1(n3754), .B2(n893), .A(n6403), .ZN(n13183) );
  oai21d1 U1685 ( .B1(n3756), .B2(n893), .A(n4751), .ZN(n13184) );
  oai21d1 U1686 ( .B1(n3758), .B2(n893), .A(n6641), .ZN(n13185) );
  oai21d1 U1687 ( .B1(n3760), .B2(n893), .A(n5298), .ZN(n13186) );
  oai21d1 U1688 ( .B1(n3762), .B2(n893), .A(n6953), .ZN(n13187) );
  oai21d1 U1689 ( .B1(n3763), .B2(n893), .A(n5776), .ZN(n13188) );
  oai21d1 U1691 ( .B1(n3765), .B2(n893), .A(n7255), .ZN(n13189) );
  oai21d1 U1695 ( .B1(n3768), .B2(n892), .A(n6140), .ZN(n13190) );
  oai21d1 U1696 ( .B1(n3709), .B2(n892), .A(n6200), .ZN(n13191) );
  oai21d1 U1697 ( .B1(n3711), .B2(n892), .A(n4222), .ZN(n13192) );
  oai21d1 U1698 ( .B1(n3713), .B2(n892), .A(n6502), .ZN(n13193) );
  oai21d1 U1699 ( .B1(n3714), .B2(n892), .A(n4974), .ZN(n13194) );
  oai21d1 U1700 ( .B1(n3716), .B2(n891), .A(n6701), .ZN(n13195) );
  oai21d1 U1701 ( .B1(n3718), .B2(n891), .A(n5459), .ZN(n13196) );
  oai21d1 U1702 ( .B1(n3720), .B2(n891), .A(n7045), .ZN(n13197) );
  oai21d1 U1703 ( .B1(n3722), .B2(n891), .A(n5862), .ZN(n13198) );
  oai21d1 U1704 ( .B1(n3724), .B2(n891), .A(n6270), .ZN(n13199) );
  oai21d1 U1705 ( .B1(n3726), .B2(n891), .A(n12172), .ZN(n13200) );
  oai21d1 U1706 ( .B1(n3727), .B2(n891), .A(n6550), .ZN(n13201) );
  oai21d1 U1707 ( .B1(n3729), .B2(n891), .A(n5110), .ZN(n13202) );
  oai21d1 U1708 ( .B1(n3731), .B2(n891), .A(n12130), .ZN(n13203) );
  oai21d1 U1709 ( .B1(n3733), .B2(n890), .A(n5585), .ZN(n13204) );
  oai21d1 U1710 ( .B1(n3735), .B2(n890), .A(n7105), .ZN(n13205) );
  oai21d1 U1711 ( .B1(n3737), .B2(n890), .A(n5959), .ZN(n13206) );
  oai21d1 U1712 ( .B1(n3739), .B2(n890), .A(n6348), .ZN(n13207) );
  oai21d1 U1713 ( .B1(n3741), .B2(n890), .A(n4512), .ZN(n13208) );
  oai21d1 U1714 ( .B1(n3743), .B2(n890), .A(n6589), .ZN(n13209) );
  oai21d1 U1715 ( .B1(n3745), .B2(n890), .A(n5205), .ZN(n13210) );
  oai21d1 U1716 ( .B1(n3747), .B2(n890), .A(n6884), .ZN(n13211) );
  oai21d1 U1717 ( .B1(n3749), .B2(n890), .A(n5704), .ZN(n13212) );
  oai21d1 U1718 ( .B1(n3750), .B2(n889), .A(n7183), .ZN(n13213) );
  oai21d1 U1719 ( .B1(n3752), .B2(n889), .A(n6070), .ZN(n13214) );
  oai21d1 U1720 ( .B1(n3754), .B2(n889), .A(n6411), .ZN(n13215) );
  oai21d1 U1721 ( .B1(n3756), .B2(n889), .A(n4754), .ZN(n13216) );
  oai21d1 U1722 ( .B1(n3758), .B2(n889), .A(n6646), .ZN(n13217) );
  oai21d1 U1723 ( .B1(n3760), .B2(n889), .A(n5312), .ZN(n13218) );
  oai21d1 U1724 ( .B1(n3762), .B2(n889), .A(n12120), .ZN(n13219) );
  oai21d1 U1725 ( .B1(n3763), .B2(n889), .A(n5782), .ZN(n13220) );
  oai21d1 U1726 ( .B1(n3765), .B2(n889), .A(n7260), .ZN(n13221) );
  oai21d1 U1731 ( .B1(n3768), .B2(n885), .A(n6146), .ZN(n13222) );
  oai21d1 U1732 ( .B1(n3709), .B2(n885), .A(n6207), .ZN(n13223) );
  oai21d1 U1734 ( .B1(n3711), .B2(n885), .A(n4292), .ZN(n13224) );
  oai21d1 U1736 ( .B1(n3713), .B2(n885), .A(n6507), .ZN(n13225) );
  oai21d1 U1738 ( .B1(n3714), .B2(n885), .A(n4976), .ZN(n13226) );
  oai21d1 U1741 ( .B1(n3716), .B2(n885), .A(n6707), .ZN(n13227) );
  oai21d1 U1743 ( .B1(n3718), .B2(n885), .A(n5466), .ZN(n13228) );
  oai21d1 U1745 ( .B1(n3720), .B2(n885), .A(n7047), .ZN(n13229) );
  oai21d1 U1747 ( .B1(n3722), .B2(n885), .A(n5864), .ZN(n13230) );
  oai21d1 U1749 ( .B1(n3724), .B2(n886), .A(n6273), .ZN(n13231) );
  oai21d1 U1751 ( .B1(n3726), .B2(n886), .A(n4342), .ZN(n13232) );
  oai21d1 U1753 ( .B1(n3727), .B2(n886), .A(n6552), .ZN(n13233) );
  oai21d1 U1755 ( .B1(n3729), .B2(n886), .A(n5113), .ZN(n13234) );
  oai21d1 U1758 ( .B1(n3731), .B2(n886), .A(n6813), .ZN(n13235) );
  oai21d1 U1760 ( .B1(n3733), .B2(n886), .A(n5591), .ZN(n13236) );
  oai21d1 U1762 ( .B1(n3735), .B2(n886), .A(n7109), .ZN(n13237) );
  oai21d1 U1765 ( .B1(n3737), .B2(n886), .A(n5964), .ZN(n13238) );
  oai21d1 U1767 ( .B1(n3739), .B2(n886), .A(n6355), .ZN(n13239) );
  oai21d1 U1769 ( .B1(n3741), .B2(n887), .A(n4608), .ZN(n13240) );
  oai21d1 U1771 ( .B1(n3743), .B2(n887), .A(n6590), .ZN(n13241) );
  oai21d1 U1773 ( .B1(n3745), .B2(n887), .A(n5220), .ZN(n13242) );
  oai21d1 U1775 ( .B1(n3747), .B2(n887), .A(n12126), .ZN(n13243) );
  oai21d1 U1777 ( .B1(n3749), .B2(n887), .A(n12164), .ZN(n13244) );
  oai21d1 U1779 ( .B1(n3750), .B2(n887), .A(n7184), .ZN(n13245) );
  oai21d1 U1783 ( .B1(n3752), .B2(n887), .A(n6072), .ZN(n13246) );
  oai21d1 U1785 ( .B1(n3754), .B2(n887), .A(n6413), .ZN(n13247) );
  oai21d1 U1788 ( .B1(n3756), .B2(n887), .A(n4871), .ZN(n13248) );
  oai21d1 U1791 ( .B1(n3758), .B2(n888), .A(n6653), .ZN(n13249) );
  oai21d1 U1794 ( .B1(n3760), .B2(n888), .A(n5315), .ZN(n13250) );
  oai21d1 U1797 ( .B1(n3762), .B2(n888), .A(n6975), .ZN(n13251) );
  oai21d1 U1800 ( .B1(n3763), .B2(n888), .A(n5785), .ZN(n13252) );
  oai21d1 U1808 ( .B1(n948), .B2(n3768), .A(n12163), .ZN(n13253) );
  oaim22d1 U1817 ( .A1(n12204), .A2(n4234), .B1(n510), .B2(n4234), .ZN(n13254)
         );
  oaim22d1 U1818 ( .A1(n12205), .A2(n4234), .B1(N3181), .B2(n4234), .ZN(n13255) );
  oaim22d1 U1819 ( .A1(n12206), .A2(n4234), .B1(N3180), .B2(n4234), .ZN(n13256) );
  oaim22d1 U1820 ( .A1(n12207), .A2(n4234), .B1(N3179), .B2(n4234), .ZN(n13257) );
  oaim22d1 U1821 ( .A1(n12208), .A2(n4234), .B1(N3976), .B2(n4234), .ZN(n13258) );
  oaim22d1 U1822 ( .A1(n12209), .A2(n4234), .B1(n955), .B2(n4234), .ZN(n13259)
         );
  oaim22d1 U1823 ( .A1(n12210), .A2(n4234), .B1(N3974), .B2(n4234), .ZN(n13260) );
  oaim22d1 U1824 ( .A1(n12211), .A2(n4234), .B1(N3973), .B2(n4234), .ZN(n13261) );
  oaim22d1 U1825 ( .A1(n12212), .A2(n4234), .B1(N3972), .B2(n4234), .ZN(n13262) );
  oai221d1 U1828 ( .B1(n2757), .B2(n12091), .C1(n12092), .C2(n4240), .A(n4241), 
        .ZN(n13263) );
  oai221d1 U1829 ( .B1(n2757), .B2(n12089), .C1(n12090), .C2(n4240), .A(n4241), 
        .ZN(n13264) );
  oai221d1 U1830 ( .B1(n2757), .B2(n12087), .C1(n12088), .C2(n4240), .A(n4241), 
        .ZN(n13265) );
  oai221d1 U1831 ( .B1(n2757), .B2(n12085), .C1(n12086), .C2(n4240), .A(n4241), 
        .ZN(n13266) );
  oai221d1 U1832 ( .B1(n2757), .B2(n12083), .C1(n12084), .C2(n4240), .A(n4241), 
        .ZN(n13267) );
  oai221d1 U1833 ( .B1(n2757), .B2(n12081), .C1(n12082), .C2(n4240), .A(n4241), 
        .ZN(n13268) );
  oai221d1 U1834 ( .B1(n2757), .B2(n12079), .C1(n12080), .C2(n4240), .A(n4241), 
        .ZN(n13269) );
  oai221d1 U1835 ( .B1(n2757), .B2(n12077), .C1(n12078), .C2(n4240), .A(n4241), 
        .ZN(n13270) );
  oai221d1 U1836 ( .B1(n2757), .B2(n12075), .C1(n12076), .C2(n4240), .A(n4241), 
        .ZN(n13271) );
  oai221d1 U1839 ( .B1(n2756), .B2(n12092), .C1(n2744), .C2(n496), .A(n4241), 
        .ZN(n13272) );
  oai221d1 U1841 ( .B1(n2756), .B2(n12090), .C1(n2745), .C2(n496), .A(n4241), 
        .ZN(n13273) );
  oai221d1 U1843 ( .B1(n2756), .B2(n12088), .C1(n2746), .C2(n496), .A(n4241), 
        .ZN(n13274) );
  oai221d1 U1845 ( .B1(n2756), .B2(n12086), .C1(n2747), .C2(n496), .A(n4241), 
        .ZN(n13275) );
  oai221d1 U1847 ( .B1(n2756), .B2(n12084), .C1(n2748), .C2(n496), .A(n4241), 
        .ZN(n13276) );
  oai221d1 U1849 ( .B1(n2756), .B2(n12082), .C1(n2749), .C2(n496), .A(n4241), 
        .ZN(n13277) );
  oai221d1 U1851 ( .B1(n2756), .B2(n12080), .C1(n2750), .C2(n496), .A(n4241), 
        .ZN(n13278) );
  oai221d1 U1853 ( .B1(n2756), .B2(n12078), .C1(n2751), .C2(n496), .A(n4241), 
        .ZN(n13279) );
  oai221d1 U1855 ( .B1(n2756), .B2(n12076), .C1(n2752), .C2(n496), .A(n4241), 
        .ZN(n13280) );
  xr02d1 U2491 ( .A1(n2778), .A2(n4375), .Z(n13793) );
  oai22d1 U2497 ( .A1(new_reference_is_done), .A2(n880), .B1(n3707), .B2(n2787), .ZN(n13794) );
  oai21d1 U2500 ( .B1(new_reference_is_done), .B2(n3657), .A(n493), .ZN(n4254)
         );
  xr02d1 U2522 ( .A1(n12468), .A2(n12724), .Z(N5019) );
  xr02d1 U2523 ( .A1(n12467), .A2(n12723), .Z(N5018) );
  xr02d1 U2524 ( .A1(n12466), .A2(n12722), .Z(N5017) );
  xr02d1 U2525 ( .A1(n12465), .A2(n12721), .Z(N5016) );
  xr02d1 U2526 ( .A1(n12464), .A2(n12720), .Z(N5015) );
  xr02d1 U2527 ( .A1(n12463), .A2(n12719), .Z(N5014) );
  xr02d1 U2528 ( .A1(n12462), .A2(n12718), .Z(N5013) );
  xr02d1 U2529 ( .A1(n12461), .A2(n12717), .Z(N5012) );
  xr02d1 U2530 ( .A1(n12460), .A2(n12716), .Z(N5011) );
  xr02d1 U2531 ( .A1(n12459), .A2(n12715), .Z(N5010) );
  xr02d1 U2532 ( .A1(n12458), .A2(n12714), .Z(N5009) );
  xr02d1 U2533 ( .A1(n12457), .A2(n12713), .Z(N5008) );
  xr02d1 U2534 ( .A1(n12456), .A2(n12712), .Z(N5007) );
  xr02d1 U2535 ( .A1(n12455), .A2(n12711), .Z(N5006) );
  xr02d1 U2536 ( .A1(n12454), .A2(n12710), .Z(N5005) );
  xr02d1 U2537 ( .A1(n12453), .A2(n12709), .Z(N5004) );
  xr02d1 U2538 ( .A1(n12452), .A2(n12708), .Z(N5003) );
  xr02d1 U2539 ( .A1(n12451), .A2(n12707), .Z(N5002) );
  xr02d1 U2540 ( .A1(n12450), .A2(n12706), .Z(N5001) );
  xr02d1 U2541 ( .A1(n12449), .A2(n12705), .Z(N5000) );
  xr02d1 U2542 ( .A1(n12448), .A2(n12704), .Z(N4999) );
  xr02d1 U2543 ( .A1(n12447), .A2(n12703), .Z(N4998) );
  xr02d1 U2544 ( .A1(n12446), .A2(n12702), .Z(N4997) );
  xr02d1 U2545 ( .A1(n12445), .A2(n12701), .Z(N4996) );
  xr02d1 U2546 ( .A1(n12444), .A2(n12700), .Z(N4995) );
  xr02d1 U2547 ( .A1(n12443), .A2(n12699), .Z(N4994) );
  xr02d1 U2548 ( .A1(n12442), .A2(n12698), .Z(N4993) );
  xr02d1 U2549 ( .A1(n12441), .A2(n12697), .Z(N4992) );
  xr02d1 U2550 ( .A1(n12440), .A2(n12696), .Z(N4991) );
  xr02d1 U2551 ( .A1(n12439), .A2(n12695), .Z(N4990) );
  xr02d1 U2552 ( .A1(n12438), .A2(n12694), .Z(N4989) );
  xr02d1 U2553 ( .A1(n12437), .A2(n12693), .Z(N4988) );
  xr02d1 U2554 ( .A1(n12436), .A2(n12692), .Z(N4987) );
  xr02d1 U2555 ( .A1(n12435), .A2(n12691), .Z(N4986) );
  xr02d1 U2556 ( .A1(n12434), .A2(n12690), .Z(N4985) );
  xr02d1 U2557 ( .A1(n12433), .A2(n12689), .Z(N4984) );
  xr02d1 U2558 ( .A1(n12432), .A2(n12688), .Z(N4983) );
  xr02d1 U2559 ( .A1(n12431), .A2(n12687), .Z(N4982) );
  xr02d1 U2560 ( .A1(n12430), .A2(n12686), .Z(N4981) );
  xr02d1 U2561 ( .A1(n12429), .A2(n12685), .Z(N4980) );
  xr02d1 U2562 ( .A1(n12428), .A2(n12684), .Z(N4979) );
  xr02d1 U2563 ( .A1(n12427), .A2(n12683), .Z(N4978) );
  xr02d1 U2564 ( .A1(n12426), .A2(n12682), .Z(N4977) );
  xr02d1 U2565 ( .A1(n12425), .A2(n12681), .Z(N4976) );
  xr02d1 U2566 ( .A1(n12424), .A2(n12680), .Z(N4975) );
  xr02d1 U2567 ( .A1(n12423), .A2(n12679), .Z(N4974) );
  xr02d1 U2568 ( .A1(n12422), .A2(n12678), .Z(N4973) );
  xr02d1 U2569 ( .A1(n12421), .A2(n12677), .Z(N4972) );
  xr02d1 U2570 ( .A1(n12420), .A2(n12676), .Z(N4971) );
  xr02d1 U2571 ( .A1(n12419), .A2(n12675), .Z(N4970) );
  xr02d1 U2572 ( .A1(n12418), .A2(n12674), .Z(N4969) );
  xr02d1 U2573 ( .A1(n12417), .A2(n12673), .Z(N4968) );
  xr02d1 U2574 ( .A1(n12416), .A2(n12672), .Z(N4967) );
  xr02d1 U2575 ( .A1(n12415), .A2(n12671), .Z(N4966) );
  xr02d1 U2576 ( .A1(n12414), .A2(n12670), .Z(N4965) );
  xr02d1 U2577 ( .A1(n12413), .A2(n12669), .Z(N4964) );
  xr02d1 U2578 ( .A1(n12412), .A2(n12668), .Z(N4963) );
  xr02d1 U2579 ( .A1(n12411), .A2(n12667), .Z(N4962) );
  xr02d1 U2580 ( .A1(n12410), .A2(n12666), .Z(N4961) );
  xr02d1 U2581 ( .A1(n12409), .A2(n12665), .Z(N4960) );
  xr02d1 U2582 ( .A1(n12408), .A2(n12664), .Z(N4959) );
  xr02d1 U2583 ( .A1(n12407), .A2(n12663), .Z(N4958) );
  xr02d1 U2584 ( .A1(n12406), .A2(n12662), .Z(N4957) );
  xr02d1 U2585 ( .A1(n12405), .A2(n12661), .Z(N4956) );
  xr02d1 U2586 ( .A1(n12404), .A2(n12660), .Z(N4955) );
  xr02d1 U2587 ( .A1(n12403), .A2(n12659), .Z(N4954) );
  xr02d1 U2588 ( .A1(n12402), .A2(n12658), .Z(N4953) );
  xr02d1 U2589 ( .A1(n12401), .A2(n12657), .Z(N4952) );
  xr02d1 U2590 ( .A1(n12400), .A2(n12656), .Z(N4951) );
  xr02d1 U2591 ( .A1(n12399), .A2(n12655), .Z(N4950) );
  xr02d1 U2592 ( .A1(n12398), .A2(n12654), .Z(N4949) );
  xr02d1 U2593 ( .A1(n12397), .A2(n12653), .Z(N4948) );
  xr02d1 U2594 ( .A1(n12396), .A2(n12652), .Z(N4947) );
  xr02d1 U2595 ( .A1(n12395), .A2(n12651), .Z(N4946) );
  xr02d1 U2596 ( .A1(n12394), .A2(n12650), .Z(N4945) );
  xr02d1 U2597 ( .A1(n12393), .A2(n12649), .Z(N4944) );
  xr02d1 U2598 ( .A1(n12392), .A2(n12648), .Z(N4943) );
  xr02d1 U2599 ( .A1(n12391), .A2(n12647), .Z(N4942) );
  xr02d1 U2600 ( .A1(n12390), .A2(n12646), .Z(N4941) );
  xr02d1 U2601 ( .A1(n12389), .A2(n12645), .Z(N4940) );
  xr02d1 U2602 ( .A1(n12388), .A2(n12644), .Z(N4939) );
  xr02d1 U2603 ( .A1(n12387), .A2(n12643), .Z(N4938) );
  xr02d1 U2604 ( .A1(n12386), .A2(n12642), .Z(N4937) );
  xr02d1 U2605 ( .A1(n12385), .A2(n12641), .Z(N4936) );
  xr02d1 U2606 ( .A1(n12384), .A2(n12640), .Z(N4935) );
  xr02d1 U2607 ( .A1(n12383), .A2(n12639), .Z(N4934) );
  xr02d1 U2608 ( .A1(n12382), .A2(n12638), .Z(N4933) );
  xr02d1 U2609 ( .A1(n12381), .A2(n12637), .Z(N4932) );
  xr02d1 U2610 ( .A1(n12380), .A2(n12636), .Z(N4931) );
  xr02d1 U2611 ( .A1(n12379), .A2(n12635), .Z(N4930) );
  xr02d1 U2612 ( .A1(n12378), .A2(n12634), .Z(N4929) );
  xr02d1 U2613 ( .A1(n12377), .A2(n12633), .Z(N4928) );
  xr02d1 U2614 ( .A1(n12376), .A2(n12632), .Z(N4927) );
  xr02d1 U2615 ( .A1(n12375), .A2(n12631), .Z(N4926) );
  xr02d1 U2616 ( .A1(n12374), .A2(n12630), .Z(N4925) );
  xr02d1 U2617 ( .A1(n12373), .A2(n12629), .Z(N4924) );
  xr02d1 U2618 ( .A1(n12372), .A2(n12628), .Z(N4923) );
  xr02d1 U2619 ( .A1(n12371), .A2(n12627), .Z(N4922) );
  xr02d1 U2620 ( .A1(n12370), .A2(n12626), .Z(N4921) );
  xr02d1 U2621 ( .A1(n12369), .A2(n12625), .Z(N4920) );
  xr02d1 U2622 ( .A1(n12368), .A2(n12624), .Z(N4919) );
  xr02d1 U2623 ( .A1(n12367), .A2(n12623), .Z(N4918) );
  xr02d1 U2624 ( .A1(n12366), .A2(n12622), .Z(N4917) );
  xr02d1 U2625 ( .A1(n12365), .A2(n12621), .Z(N4916) );
  xr02d1 U2626 ( .A1(n12364), .A2(n12620), .Z(N4915) );
  xr02d1 U2627 ( .A1(n12363), .A2(n12619), .Z(N4914) );
  xr02d1 U2628 ( .A1(n12362), .A2(n12618), .Z(N4913) );
  xr02d1 U2629 ( .A1(n12361), .A2(n12617), .Z(N4912) );
  xr02d1 U2630 ( .A1(n12360), .A2(n12616), .Z(N4911) );
  xr02d1 U2631 ( .A1(n12359), .A2(n12615), .Z(N4910) );
  xr02d1 U2632 ( .A1(n12358), .A2(n12614), .Z(N4909) );
  xr02d1 U2633 ( .A1(n12357), .A2(n12613), .Z(N4908) );
  xr02d1 U2634 ( .A1(n12356), .A2(n12612), .Z(N4907) );
  xr02d1 U2635 ( .A1(n12355), .A2(n12611), .Z(N4906) );
  xr02d1 U2636 ( .A1(n12354), .A2(n12610), .Z(N4905) );
  xr02d1 U2637 ( .A1(n12353), .A2(n12609), .Z(N4904) );
  xr02d1 U2638 ( .A1(n12352), .A2(n12608), .Z(N4903) );
  xr02d1 U2639 ( .A1(n12351), .A2(n12607), .Z(N4902) );
  xr02d1 U2640 ( .A1(n12350), .A2(n12606), .Z(N4901) );
  xr02d1 U2641 ( .A1(n12349), .A2(n12605), .Z(N4900) );
  xr02d1 U2642 ( .A1(n12348), .A2(n12604), .Z(N4899) );
  xr02d1 U2643 ( .A1(n12347), .A2(n12603), .Z(N4898) );
  xr02d1 U2644 ( .A1(n12346), .A2(n12602), .Z(N4897) );
  xr02d1 U2645 ( .A1(n12345), .A2(n12601), .Z(N4896) );
  xr02d1 U2646 ( .A1(n12344), .A2(n12600), .Z(N4895) );
  xr02d1 U2647 ( .A1(n12343), .A2(n12599), .Z(N4894) );
  xr02d1 U2648 ( .A1(n12342), .A2(n12598), .Z(N4893) );
  xr02d1 U2649 ( .A1(n12341), .A2(n12597), .Z(N4892) );
  xr02d1 U2650 ( .A1(n12340), .A2(n12596), .Z(N4891) );
  xr02d1 U2651 ( .A1(n12339), .A2(n12595), .Z(N4890) );
  xr02d1 U2652 ( .A1(n12338), .A2(n12594), .Z(N4889) );
  xr02d1 U2653 ( .A1(n12337), .A2(n12593), .Z(N4888) );
  xr02d1 U2654 ( .A1(n12336), .A2(n12592), .Z(N4887) );
  xr02d1 U2655 ( .A1(n12335), .A2(n12591), .Z(N4886) );
  xr02d1 U2656 ( .A1(n12334), .A2(n12590), .Z(N4885) );
  xr02d1 U2657 ( .A1(n12333), .A2(n12589), .Z(N4884) );
  xr02d1 U2658 ( .A1(n12332), .A2(n12588), .Z(N4883) );
  xr02d1 U2659 ( .A1(n12331), .A2(n12587), .Z(N4882) );
  xr02d1 U2660 ( .A1(n12330), .A2(n12586), .Z(N4881) );
  xr02d1 U2661 ( .A1(n12329), .A2(n12585), .Z(N4880) );
  xr02d1 U2662 ( .A1(n12328), .A2(n12584), .Z(N4879) );
  xr02d1 U2663 ( .A1(n12327), .A2(n12583), .Z(N4878) );
  xr02d1 U2664 ( .A1(n12326), .A2(n12582), .Z(N4877) );
  xr02d1 U2665 ( .A1(n12325), .A2(n12581), .Z(N4876) );
  xr02d1 U2666 ( .A1(n12324), .A2(n12580), .Z(N4875) );
  xr02d1 U2667 ( .A1(n12323), .A2(n12579), .Z(N4874) );
  xr02d1 U2668 ( .A1(n12322), .A2(n12578), .Z(N4873) );
  xr02d1 U2669 ( .A1(n12321), .A2(n12577), .Z(N4872) );
  xr02d1 U2670 ( .A1(n12320), .A2(n12576), .Z(N4871) );
  xr02d1 U2671 ( .A1(n12319), .A2(n12575), .Z(N4870) );
  xr02d1 U2672 ( .A1(n12318), .A2(n12574), .Z(N4869) );
  xr02d1 U2673 ( .A1(n12317), .A2(n12573), .Z(N4868) );
  xr02d1 U2674 ( .A1(n12316), .A2(n12572), .Z(N4867) );
  xr02d1 U2675 ( .A1(n12315), .A2(n12571), .Z(N4866) );
  xr02d1 U2676 ( .A1(n12314), .A2(n12570), .Z(N4865) );
  xr02d1 U2677 ( .A1(n12313), .A2(n12569), .Z(N4864) );
  xr02d1 U2678 ( .A1(n12312), .A2(n12568), .Z(N4863) );
  xr02d1 U2679 ( .A1(n12311), .A2(n12567), .Z(N4862) );
  xr02d1 U2680 ( .A1(n12310), .A2(n12566), .Z(N4861) );
  xr02d1 U2681 ( .A1(n12309), .A2(n12565), .Z(N4860) );
  xr02d1 U2682 ( .A1(n12308), .A2(n12564), .Z(N4859) );
  xr02d1 U2683 ( .A1(n12307), .A2(n12563), .Z(N4858) );
  xr02d1 U2684 ( .A1(n12306), .A2(n12562), .Z(N4857) );
  xr02d1 U2685 ( .A1(n12305), .A2(n12561), .Z(N4856) );
  xr02d1 U2686 ( .A1(n12304), .A2(n12560), .Z(N4855) );
  xr02d1 U2687 ( .A1(n12303), .A2(n12559), .Z(N4854) );
  xr02d1 U2688 ( .A1(n12302), .A2(n12558), .Z(N4853) );
  xr02d1 U2689 ( .A1(n12301), .A2(n12557), .Z(N4852) );
  xr02d1 U2690 ( .A1(n12300), .A2(n12556), .Z(N4851) );
  xr02d1 U2691 ( .A1(n12299), .A2(n12555), .Z(N4850) );
  xr02d1 U2692 ( .A1(n12298), .A2(n12554), .Z(N4849) );
  xr02d1 U2693 ( .A1(n12297), .A2(n12553), .Z(N4848) );
  xr02d1 U2694 ( .A1(n12296), .A2(n12552), .Z(N4847) );
  xr02d1 U2695 ( .A1(n12295), .A2(n12551), .Z(N4846) );
  xr02d1 U2696 ( .A1(n12294), .A2(n12550), .Z(N4845) );
  xr02d1 U2697 ( .A1(n12293), .A2(n12549), .Z(N4844) );
  xr02d1 U2698 ( .A1(n12292), .A2(n12548), .Z(N4843) );
  xr02d1 U2699 ( .A1(n12291), .A2(n12547), .Z(N4842) );
  xr02d1 U2700 ( .A1(n12290), .A2(n12546), .Z(N4841) );
  xr02d1 U2701 ( .A1(n12289), .A2(n12545), .Z(N4840) );
  xr02d1 U2702 ( .A1(n12288), .A2(n12544), .Z(N4839) );
  xr02d1 U2703 ( .A1(n12287), .A2(n12543), .Z(N4838) );
  xr02d1 U2704 ( .A1(n12286), .A2(n12542), .Z(N4837) );
  xr02d1 U2705 ( .A1(n12285), .A2(n12541), .Z(N4836) );
  xr02d1 U2706 ( .A1(n12284), .A2(n12540), .Z(N4835) );
  xr02d1 U2707 ( .A1(n12283), .A2(n12539), .Z(N4834) );
  xr02d1 U2708 ( .A1(n12282), .A2(n12538), .Z(N4833) );
  xr02d1 U2709 ( .A1(n12281), .A2(n12537), .Z(N4832) );
  xr02d1 U2710 ( .A1(n12280), .A2(n12536), .Z(N4831) );
  xr02d1 U2711 ( .A1(n12279), .A2(n12535), .Z(N4830) );
  xr02d1 U2712 ( .A1(n12278), .A2(n12534), .Z(N4829) );
  xr02d1 U2713 ( .A1(n12277), .A2(n12533), .Z(N4828) );
  xr02d1 U2714 ( .A1(n12276), .A2(n12532), .Z(N4827) );
  xr02d1 U2715 ( .A1(n12275), .A2(n12531), .Z(N4826) );
  xr02d1 U2716 ( .A1(n12274), .A2(n12530), .Z(N4825) );
  xr02d1 U2717 ( .A1(n12273), .A2(n12529), .Z(N4824) );
  xr02d1 U2718 ( .A1(n12272), .A2(n12528), .Z(N4823) );
  xr02d1 U2719 ( .A1(n12271), .A2(n12527), .Z(N4822) );
  xr02d1 U2720 ( .A1(n12270), .A2(n12526), .Z(N4821) );
  xr02d1 U2721 ( .A1(n12269), .A2(n12525), .Z(N4820) );
  xr02d1 U2722 ( .A1(n12268), .A2(n12524), .Z(N4819) );
  xr02d1 U2723 ( .A1(n12267), .A2(n12523), .Z(N4818) );
  xr02d1 U2724 ( .A1(n12266), .A2(n12522), .Z(N4817) );
  xr02d1 U2725 ( .A1(n12265), .A2(n12521), .Z(N4816) );
  xr02d1 U2726 ( .A1(n12264), .A2(n12520), .Z(N4815) );
  xr02d1 U2727 ( .A1(n12263), .A2(n12519), .Z(N4814) );
  xr02d1 U2728 ( .A1(n12262), .A2(n12518), .Z(N4813) );
  xr02d1 U2729 ( .A1(n12261), .A2(n12517), .Z(N4812) );
  xr02d1 U2730 ( .A1(n12260), .A2(n12516), .Z(N4811) );
  xr02d1 U2731 ( .A1(n12259), .A2(n12515), .Z(N4810) );
  xr02d1 U2732 ( .A1(n12258), .A2(n12514), .Z(N4809) );
  xr02d1 U2733 ( .A1(n12257), .A2(n12513), .Z(N4808) );
  xr02d1 U2734 ( .A1(n12256), .A2(n12512), .Z(N4807) );
  xr02d1 U2735 ( .A1(n12255), .A2(n12511), .Z(N4806) );
  xr02d1 U2736 ( .A1(n12254), .A2(n12510), .Z(N4805) );
  xr02d1 U2737 ( .A1(n12253), .A2(n12509), .Z(N4804) );
  xr02d1 U2738 ( .A1(n12252), .A2(n12508), .Z(N4803) );
  xr02d1 U2739 ( .A1(n12251), .A2(n12507), .Z(N4802) );
  xr02d1 U2740 ( .A1(n12250), .A2(n12506), .Z(N4801) );
  xr02d1 U2741 ( .A1(n12249), .A2(n12505), .Z(N4800) );
  xr02d1 U2742 ( .A1(n12248), .A2(n12504), .Z(N4799) );
  xr02d1 U2743 ( .A1(n12247), .A2(n12503), .Z(N4798) );
  xr02d1 U2744 ( .A1(n12246), .A2(n12502), .Z(N4797) );
  xr02d1 U2745 ( .A1(n12245), .A2(n12501), .Z(N4796) );
  xr02d1 U2746 ( .A1(n12244), .A2(n12500), .Z(N4795) );
  xr02d1 U2747 ( .A1(n12243), .A2(n12499), .Z(N4794) );
  xr02d1 U2748 ( .A1(n12242), .A2(n12498), .Z(N4793) );
  xr02d1 U2749 ( .A1(n12241), .A2(n12497), .Z(N4792) );
  xr02d1 U2750 ( .A1(n12240), .A2(n12496), .Z(N4791) );
  xr02d1 U2751 ( .A1(n12239), .A2(n12495), .Z(N4790) );
  xr02d1 U2752 ( .A1(n12238), .A2(n12494), .Z(N4789) );
  xr02d1 U2753 ( .A1(n12237), .A2(n12493), .Z(N4788) );
  xr02d1 U2754 ( .A1(n12236), .A2(n12492), .Z(N4787) );
  xr02d1 U2755 ( .A1(n12235), .A2(n12491), .Z(N4786) );
  xr02d1 U2756 ( .A1(n12234), .A2(n12490), .Z(N4785) );
  xr02d1 U2757 ( .A1(n12233), .A2(n12489), .Z(N4784) );
  xr02d1 U2758 ( .A1(n12232), .A2(n12488), .Z(N4783) );
  xr02d1 U2759 ( .A1(n12231), .A2(n12487), .Z(N4782) );
  xr02d1 U2760 ( .A1(n12230), .A2(n12486), .Z(N4781) );
  xr02d1 U2761 ( .A1(n12229), .A2(n12485), .Z(N4780) );
  xr02d1 U2762 ( .A1(n12228), .A2(n12484), .Z(N4779) );
  xr02d1 U2763 ( .A1(n12227), .A2(n12483), .Z(N4778) );
  xr02d1 U2764 ( .A1(n12226), .A2(n12482), .Z(N4777) );
  xr02d1 U2765 ( .A1(n12225), .A2(n12481), .Z(N4776) );
  xr02d1 U2766 ( .A1(n12224), .A2(n12480), .Z(N4775) );
  xr02d1 U2767 ( .A1(n12223), .A2(n12479), .Z(N4774) );
  xr02d1 U2768 ( .A1(n12222), .A2(n12478), .Z(N4773) );
  xr02d1 U2769 ( .A1(n12221), .A2(n12477), .Z(N4772) );
  xr02d1 U2770 ( .A1(n12220), .A2(n12476), .Z(N4771) );
  xr02d1 U2771 ( .A1(n12219), .A2(n12475), .Z(N4770) );
  xr02d1 U2772 ( .A1(n12218), .A2(n12474), .Z(N4769) );
  xr02d1 U2773 ( .A1(n12217), .A2(n12473), .Z(N4768) );
  xr02d1 U2774 ( .A1(n12216), .A2(n12472), .Z(N4767) );
  xr02d1 U2775 ( .A1(n12215), .A2(n12471), .Z(N4766) );
  xr02d1 U2776 ( .A1(n12214), .A2(n12470), .Z(N4765) );
  xr02d1 U2777 ( .A1(n12213), .A2(n12469), .Z(N4764) );
  oai311d1 U2807 ( .C1(n7240), .C2(n4434), .C3(n4435), .A(n3784), .B(n3773), 
        .ZN(n4430) );
  aoi321d1 U2808 ( .C1(n3528), .C2(n4683), .C3(n4440), .B1(n3568), .B2(n4442), 
        .A(n4443), .ZN(n4434) );
  aon211d1 U2810 ( .C1(n4447), .C2(n4448), .B(n4449), .A(n4681), .ZN(n4445) );
  aoi21d1 U2811 ( .B1(n3535), .B2(n4452), .A(n4453), .ZN(n4448) );
  aoi31d1 U2812 ( .B1(n4454), .B2(n4681), .B3(n4455), .A(n4456), .ZN(n4453) );
  aoi31d1 U2813 ( .B1(n3561), .B2(n4458), .B3(n3537), .A(n4460), .ZN(n4455) );
  aoi311d1 U2814 ( .C1(n4461), .C2(n4441), .C3(n4463), .A(n3541), .B(n4465), 
        .ZN(n4460) );
  aoi22d1 U2815 ( .A1(n4466), .A2(n4467), .B1(n4468), .B2(n4469), .ZN(n4463)
         );
  oai211d1 U2816 ( .C1(n4310), .C2(n3551), .A(n4472), .B(n4473), .ZN(n4469) );
  oai31d1 U2817 ( .B1(n4474), .B2(n4467), .B3(n4475), .A(n4476), .ZN(n4472) );
  oai22d1 U2818 ( .A1(n4477), .A2(n4478), .B1(n4479), .B2(n4480), .ZN(n4474)
         );
  aon211d1 U2819 ( .C1(n3473), .C2(n4482), .B(n4483), .A(n4484), .ZN(n4480) );
  oai31d1 U2821 ( .B1(n4488), .B2(n4489), .B3(n4490), .A(n3428), .ZN(n4487) );
  aoi31d1 U2822 ( .B1(n4492), .B2(n3502), .B3(n4494), .A(n4495), .ZN(n4489) );
  aoi22d1 U2823 ( .A1(n4496), .A2(n3433), .B1(n4498), .B2(n4499), .ZN(n4494)
         );
  aoi21d1 U2824 ( .B1(n4500), .B2(n4501), .A(n4502), .ZN(n4496) );
  aon211d1 U2825 ( .C1(n3435), .C2(n4504), .B(n4505), .A(n3434), .ZN(n4501) );
  oai211d1 U2826 ( .C1(n4507), .C2(n4508), .A(n4500), .B(n4509), .ZN(n4504) );
  aoi31d1 U2827 ( .B1(n3451), .B2(n4511), .B3(n3447), .A(n4513), .ZN(n4507) );
  oai211d1 U2829 ( .C1(n4516), .C2(n4517), .A(n3500), .B(n4518), .ZN(n4511) );
  aoi311d1 U2831 ( .C1(n4520), .C2(n4521), .C3(n4522), .A(n3361), .B(n3501), 
        .ZN(n4516) );
  or04d0 U2833 ( .A1(n4526), .A2(n3501), .A3(n4527), .A4(n4528), .Z(n4521) );
  aon211d1 U2835 ( .C1(n3350), .C2(n4531), .B(n4532), .A(n4528), .ZN(n4520) );
  aoi311d1 U2837 ( .C1(n4537), .C2(n4538), .C3(n3350), .A(n4539), .B(n4540), 
        .ZN(n4533) );
  oai22d1 U2839 ( .A1(n4544), .A2(n4545), .B1(n4546), .B2(n4547), .ZN(n4542)
         );
  aoi321d1 U2840 ( .C1(n4548), .C2(n3406), .C3(n4550), .B1(n3369), .B2(n3349), 
        .A(n4553), .ZN(n4544) );
  or02d0 U2841 ( .A1(n4554), .A2(n4541), .Z(n4553) );
  aoi22d1 U2843 ( .A1(n4555), .A2(n4556), .B1(n4557), .B2(n4558), .ZN(n4550)
         );
  aoi221d1 U2844 ( .B1(n4559), .B2(n4560), .C1(n3379), .C2(n4562), .A(n4563), 
        .ZN(n4556) );
  oai211d1 U2845 ( .C1(n4564), .C2(n4565), .A(n4566), .B(n4567), .ZN(n4560) );
  aoi21d1 U2846 ( .B1(n3381), .B2(n4569), .A(n4562), .ZN(n4567) );
  aoi31d1 U2848 ( .B1(n4573), .B2(n4574), .B3(n3251), .A(n3386), .ZN(n4571) );
  aor31d1 U2849 ( .B1(n4577), .B2(n4573), .B3(n4578), .A(n4579), .Z(n4574) );
  aoi22d1 U2850 ( .A1(n3273), .A2(n4581), .B1(n4582), .B2(n4583), .ZN(n4578)
         );
  aon211d1 U2851 ( .C1(n4584), .C2(n4585), .B(n4586), .A(n3327), .ZN(n4583) );
  oai22d1 U2852 ( .A1(n4588), .A2(n4589), .B1(n3320), .B2(n4591), .ZN(n4584)
         );
  aoi22d1 U2853 ( .A1(n4592), .A2(n4593), .B1(n4594), .B2(n3317), .ZN(n4588)
         );
  oai22d1 U2854 ( .A1(n4596), .A2(n4597), .B1(n4598), .B2(n4599), .ZN(n4593)
         );
  aoim31d1 U2855 ( .B1(n4600), .B2(n4601), .B3(n4602), .A(n4603), .ZN(n4596)
         );
  oan211d1 U2856 ( .C1(n5146), .C2(n4600), .B(n3279), .A(n4605), .ZN(n4603) );
  oai22d1 U2857 ( .A1(n4606), .A2(n4607), .B1(n3280), .B2(n4601), .ZN(n4600)
         );
  oai222d1 U2859 ( .A1(n4612), .A2(n4613), .B1(n4614), .B2(n4615), .C1(n4616), 
        .C2(n4617), .ZN(n4609) );
  aoi21d1 U2860 ( .B1(n4618), .B2(n3290), .A(n4620), .ZN(n4614) );
  aoi31d1 U2861 ( .B1(n4621), .B2(n4612), .B3(n4622), .A(n4623), .ZN(n4618) );
  aoi21d1 U2862 ( .B1(n4624), .B2(n4625), .A(n4626), .ZN(n4622) );
  aoi31d1 U2863 ( .B1(n4627), .B2(n3252), .B3(n4629), .A(n4630), .ZN(n4626) );
  aoi222d1 U2864 ( .A1(n4631), .A2(n4632), .B1(n3299), .B2(n4634), .C1(n3164), 
        .C2(n4636), .ZN(n4629) );
  oai211d1 U2865 ( .C1(n4637), .C2(n4638), .A(n4639), .B(n3247), .ZN(n4636) );
  aoi31d1 U2867 ( .B1(n4645), .B2(n3160), .B3(n4647), .A(n4648), .ZN(n4643) );
  aoi211d1 U2868 ( .C1(n3175), .C2(n4650), .A(n4651), .B(n4652), .ZN(n4647) );
  aoi31d1 U2869 ( .B1(n3159), .B2(images_bus[391]), .B3(n4654), .A(n4655), 
        .ZN(n4651) );
  aoi211d1 U2870 ( .C1(n3243), .C2(n4657), .A(n4658), .B(n4659), .ZN(n4654) );
  aoi31d1 U2871 ( .B1(n4660), .B2(n4661), .B3(n4662), .A(n3242), .ZN(n4658) );
  aoi21d1 U2872 ( .B1(n4664), .B2(n4665), .A(n4657), .ZN(n4662) );
  oai211d1 U2873 ( .C1(n4666), .C2(n4667), .A(n3190), .B(n4669), .ZN(n4665) );
  aoi211d1 U2874 ( .C1(n4670), .C2(n4671), .A(n4672), .B(n4673), .ZN(n4666) );
  oai22d1 U2875 ( .A1(n4674), .A2(n3194), .B1(n4676), .B2(n3197), .ZN(n4672)
         );
  aoi221d1 U2876 ( .B1(n4678), .B2(n4679), .C1(n4680), .C2(n3157), .A(n4682), 
        .ZN(n4676) );
  oai211d1 U2878 ( .C1(n3231), .C2(n4684), .A(n4685), .B(n4686), .ZN(n4679) );
  aoi221d1 U2879 ( .B1(n4687), .B2(n4688), .C1(n3215), .C2(n4690), .A(n3230), 
        .ZN(n4686) );
  oai211d1 U2880 ( .C1(n3227), .C2(n3158), .A(n4694), .B(n4695), .ZN(n4690) );
  aoi221d1 U2881 ( .B1(n4696), .B2(n4697), .C1(n3028), .C2(n4699), .A(n4700), 
        .ZN(n4695) );
  oan211d1 U2882 ( .C1(n4701), .C2(n4702), .B(n3033), .A(n4704), .ZN(n4700) );
  oai211d1 U2884 ( .C1(n4706), .C2(n4707), .A(n4708), .B(n4709), .ZN(n4699) );
  aoi22d1 U2885 ( .A1(n4710), .A2(n3021), .B1(n4712), .B2(n4713), .ZN(n4709)
         );
  aoi211d1 U2887 ( .C1(n4715), .C2(n4716), .A(n4717), .B(n4718), .ZN(n4706) );
  oai22d1 U2888 ( .A1(n3022), .A2(n4720), .B1(n4721), .B2(n4714), .ZN(n4717)
         );
  oai211d1 U2890 ( .C1(n4723), .C2(n4724), .A(n3053), .B(n4726), .ZN(n4716) );
  aoi22d1 U2891 ( .A1(n3056), .A2(n4728), .B1(n4729), .B2(n4722), .ZN(n4726)
         );
  oai221d1 U2892 ( .B1(n4730), .B2(n4731), .C1(n4732), .C2(n4733), .A(n4734), 
        .ZN(n4728) );
  aoim211d1 U2893 ( .C1(n4723), .C2(n3065), .A(n4736), .B(n4737), .ZN(n4732)
         );
  oaim22d1 U2894 ( .A1(n4738), .A2(n4739), .B1(n4740), .B2(n4741), .ZN(n4736)
         );
  aoi22d1 U2895 ( .A1(n3072), .A2(n4743), .B1(n4740), .B2(n4744), .ZN(n4738)
         );
  oai211d1 U2896 ( .C1(n3023), .C2(n3120), .A(n3080), .B(n4748), .ZN(n4743) );
  aoi22d1 U2897 ( .A1(n4749), .A2(n4750), .B1(n3117), .B2(n4752), .ZN(n4748)
         );
  oai22d1 U2898 ( .A1(n4753), .A2(n3086), .B1(n4755), .B2(n4756), .ZN(n4752)
         );
  aoi211d1 U2899 ( .C1(n4750), .C2(n4757), .A(n4758), .B(n4759), .ZN(n4755) );
  oai22d1 U2900 ( .A1(n4760), .A2(n4761), .B1(n4762), .B2(n4763), .ZN(n4758)
         );
  aoi321d1 U2901 ( .C1(n4764), .C2(n4765), .C3(n3096), .B1(n3100), .B2(n4768), 
        .A(n4769), .ZN(n4762) );
  oai21d1 U2902 ( .B1(n4760), .B2(n4770), .A(n3098), .ZN(n4769) );
  oai211d1 U2904 ( .C1(n4773), .C2(n4774), .A(n4775), .B(n2919), .ZN(n4768) );
  oai21d1 U2905 ( .B1(n4777), .B2(n4778), .A(n4765), .ZN(n4775) );
  aoi211d1 U2906 ( .C1(n4765), .C2(n4779), .A(n4780), .B(n4781), .ZN(n4773) );
  oai22d1 U2907 ( .A1(n4782), .A2(n4783), .B1(n4784), .B2(n4785), .ZN(n4780)
         );
  aoi221d1 U2908 ( .B1(n4786), .B2(n4787), .C1(n4788), .C2(n2930), .A(n4790), 
        .ZN(n4782) );
  oai321d1 U2909 ( .C1(n4791), .C2(n4792), .C3(n2933), .B1(n4794), .B2(n4795), 
        .A(n4796), .ZN(n4787) );
  aoi21d1 U2910 ( .B1(n4791), .B2(n2930), .A(n4797), .ZN(n4796) );
  aoi221d1 U2912 ( .B1(n4798), .B2(n4799), .C1(n4800), .C2(n4801), .A(n4802), 
        .ZN(n4794) );
  oai321d1 U2913 ( .C1(n4803), .C2(n4804), .C3(n4805), .B1(n4806), .B2(n4807), 
        .A(n4808), .ZN(n4799) );
  aoi21d1 U2914 ( .B1(n4801), .B2(n4803), .A(n4809), .ZN(n4808) );
  aoi211d1 U2915 ( .C1(n4810), .C2(n4811), .A(n4812), .B(n4813), .ZN(n4806) );
  aoi21d1 U2916 ( .B1(n4814), .B2(n4815), .A(n4805), .ZN(n4813) );
  oai211d1 U2917 ( .C1(n2998), .C2(n4805), .A(n4817), .B(n4818), .ZN(n4811) );
  aoi322d1 U2918 ( .C1(n2990), .C2(n4820), .C3(n4821), .A1(n4822), .A2(n4823), 
        .B1(n4824), .B2(n4825), .ZN(n4818) );
  oai211d1 U2919 ( .C1(n4826), .C2(n2932), .A(n4828), .B(n4829), .ZN(n4825) );
  aoi211d1 U2920 ( .C1(n4830), .C2(n4831), .A(n2987), .B(n4833), .ZN(n4829) );
  oan211d1 U2921 ( .C1(n4834), .C2(n2969), .B(n4836), .A(n4837), .ZN(n4833) );
  oai21d1 U2922 ( .B1(n4838), .B2(n4839), .A(n4831), .ZN(n4836) );
  aoi211d1 U2923 ( .C1(n4831), .C2(n4840), .A(n4841), .B(n4842), .ZN(n4834) );
  oai222d1 U2924 ( .A1(n4843), .A2(n2981), .B1(n4845), .B2(n4846), .C1(n2931), 
        .C2(n4848), .ZN(n4841) );
  aoi211d1 U2925 ( .C1(n4849), .C2(n4850), .A(n4851), .B(n4852), .ZN(n4845) );
  oai222d1 U2926 ( .A1(n4853), .A2(n2827), .B1(n4855), .B2(n4856), .C1(n4853), 
        .C2(n4857), .ZN(n4851) );
  aoi22d1 U2927 ( .A1(n2850), .A2(n4859), .B1(n4860), .B2(n4861), .ZN(n4855)
         );
  oai211d1 U2928 ( .C1(n4862), .C2(n4863), .A(n4864), .B(n4865), .ZN(n4859) );
  aoi21d1 U2929 ( .B1(n2855), .B2(n4867), .A(n4868), .ZN(n4865) );
  aoi21d1 U2930 ( .B1(n4869), .B2(n4870), .A(n2841), .ZN(n4868) );
  aoi211d1 U2931 ( .C1(n4872), .C2(n4867), .A(n4873), .B(n4874), .ZN(n4862) );
  oaim22d1 U2932 ( .A1(n4875), .A2(n4876), .B1(n4877), .B2(n4878), .ZN(n4873)
         );
  aoi211d1 U2933 ( .C1(n4879), .C2(n4877), .A(n4880), .B(n2873), .ZN(n4875) );
  aon211d1 U2934 ( .C1(n4882), .C2(n4883), .B(n4884), .A(n4885), .ZN(n4880) );
  aoi22d1 U2935 ( .A1(n2884), .A2(n4887), .B1(n4888), .B2(n2839), .ZN(n4883)
         );
  oai211d1 U2936 ( .C1(n2840), .C2(n4891), .A(n4892), .B(n4893), .ZN(n4887) );
  aoi22d1 U2937 ( .A1(n2907), .A2(n2839), .B1(n2905), .B2(n4896), .ZN(n4893)
         );
  aoi31d1 U2939 ( .B1(n4898), .B2(n4899), .B3(n2903), .A(n2890), .ZN(n4892) );
  oai321d1 U2940 ( .C1(n2895), .C2(n4903), .C3(n4904), .B1(n4905), .B2(n4906), 
        .A(n4907), .ZN(n4899) );
  aoi21d1 U2941 ( .B1(n4908), .B2(n4896), .A(n4909), .ZN(n4907) );
  aoim211d1 U2942 ( .C1(n4903), .C2(n4910), .A(n4911), .B(n4912), .ZN(n4905)
         );
  aoi31d1 U2943 ( .B1(n4889), .B2(n4903), .B3(n4914), .A(n2898), .ZN(n4912) );
  aoi21d1 U2948 ( .B1(n4918), .B2(n4920), .A(n4921), .ZN(n4882) );
  nd13d1 U2949 ( .A1(n4877), .A2(n4396), .A3(n4923), .ZN(n4918) );
  oai21d1 U2956 ( .B1(n4929), .B2(n4930), .A(n4931), .ZN(n4928) );
  aoim21d1 U2959 ( .B1(n4934), .B2(n2931), .A(n4935), .ZN(n4843) );
  oai21d1 U3019 ( .B1(n4997), .B2(n4490), .A(n3472), .ZN(n4486) );
  aoi211d1 U3029 ( .C1(images_bus[128]), .C2(n5009), .A(n5008), .B(n4432), 
        .ZN(N26365) );
  or04d0 U3032 ( .A1(n5018), .A2(n5019), .A3(n5020), .A4(n5021), .Z(n5014) );
  oai321d1 U3041 ( .C1(n4005), .C2(n5047), .C3(n5048), .B1(n4055), .B2(n5050), 
        .A(n5051), .ZN(n5045) );
  aoi21d1 U3042 ( .B1(n4006), .B2(n5053), .A(n5054), .ZN(n5051) );
  aoim211d1 U3043 ( .C1(n5055), .C2(images_bus[135]), .A(n5056), .B(n5057), 
        .ZN(n5047) );
  aoi21d1 U3044 ( .B1(n5058), .B2(n5059), .A(n5007), .ZN(n5057) );
  aon211d1 U3045 ( .C1(n4020), .C2(n2806), .B(n5062), .A(n4015), .ZN(n5059) );
  aoim211d1 U3047 ( .C1(n5065), .C2(n5066), .A(n5062), .B(n5067), .ZN(n5064)
         );
  aoi321d1 U3048 ( .C1(n4025), .C2(n5069), .C3(n5070), .B1(n4022), .B2(n5072), 
        .A(n5073), .ZN(n5065) );
  oai21d1 U3049 ( .B1(images_bus[141]), .B2(n5074), .A(n5075), .ZN(n5073) );
  oai211d1 U3050 ( .C1(images_bus[143]), .C2(n5076), .A(n5077), .B(n5078), 
        .ZN(n5069) );
  aoi22d1 U3051 ( .A1(n4026), .A2(n5080), .B1(n5081), .B2(n5573), .ZN(n5078)
         );
  aon211d1 U3052 ( .C1(n5082), .C2(n5083), .B(n5084), .A(n5085), .ZN(n5080) );
  aor31d1 U3053 ( .B1(n5085), .B2(n5082), .B3(n5086), .A(n5087), .Z(n5083) );
  aoi211d1 U3054 ( .C1(n5088), .C2(n5089), .A(n5090), .B(n5091), .ZN(n5086) );
  aoi31d1 U3055 ( .B1(n5092), .B2(n4481), .B3(n5094), .A(n5095), .ZN(n5091) );
  aoi22d1 U3056 ( .A1(n4036), .A2(n5097), .B1(n4046), .B2(n5099), .ZN(n5094)
         );
  aon211d1 U3057 ( .C1(n5100), .C2(n4041), .B(n5102), .A(images_bus[152]), 
        .ZN(n5097) );
  aoi22d1 U3059 ( .A1(n4038), .A2(n5105), .B1(n4042), .B2(n5107), .ZN(n5100)
         );
  oai21d1 U3060 ( .B1(n5108), .B2(n5109), .A(n4962), .ZN(n5105) );
  oai22d1 U3062 ( .A1(n5114), .A2(n5115), .B1(n5116), .B2(n5117), .ZN(n5111)
         );
  aoi221d1 U3063 ( .B1(n3912), .B2(n5119), .C1(n5120), .C2(n5121), .A(n7244), 
        .ZN(n5116) );
  oai211d1 U3064 ( .C1(n5122), .C2(n5123), .A(n5763), .B(n5114), .ZN(n5119) );
  oan211d1 U3065 ( .C1(n5125), .C2(n5278), .B(n3914), .A(n5127), .ZN(n5122) );
  aoi31d1 U3066 ( .B1(n5128), .B2(n3973), .B3(n5130), .A(n5131), .ZN(n5125) );
  aoim31d1 U3067 ( .B1(n6395), .B2(n5132), .B3(n5133), .A(n5134), .ZN(n5130)
         );
  oan211d1 U3068 ( .C1(images_bus[167]), .C2(n5135), .B(n3972), .A(n5137), 
        .ZN(n5134) );
  oai21d1 U3069 ( .B1(n5138), .B2(n5139), .A(n3964), .ZN(n5133) );
  aoi31d1 U3070 ( .B1(n5141), .B2(n6045), .B3(n5143), .A(n5144), .ZN(n5138) );
  aoi321d1 U3071 ( .C1(n3928), .C2(n3927), .C3(n5147), .B1(n3927), .B2(n5148), 
        .A(n5149), .ZN(n5143) );
  aoi31d1 U3072 ( .B1(n5150), .B2(n5151), .B3(n5192), .A(n5153), .ZN(n5147) );
  oai311d1 U3073 ( .C1(n5154), .C2(n5148), .C3(n5155), .A(n3933), .B(n5157), 
        .ZN(n5150) );
  oai211d1 U3074 ( .C1(images_bus[177]), .C2(n5158), .A(n5159), .B(n5192), 
        .ZN(n5154) );
  aon211d1 U3075 ( .C1(n5160), .C2(n5161), .B(n5162), .A(n5163), .ZN(n5159) );
  aoi31d1 U3076 ( .B1(n3941), .B2(n3971), .B3(n5166), .A(n5167), .ZN(n5160) );
  aoi221d1 U3077 ( .B1(n3939), .B2(n5169), .C1(n5170), .C2(n5171), .A(n5172), 
        .ZN(n5166) );
  oai211d1 U3078 ( .C1(images_bus[183]), .C2(n3946), .A(n5174), .B(n5175), 
        .ZN(n5171) );
  oai211d1 U3080 ( .C1(n5179), .C2(n5180), .A(n5181), .B(n3970), .ZN(n5176) );
  aoi211d1 U3082 ( .C1(n3955), .C2(n5183), .A(n5184), .B(n5185), .ZN(n5179) );
  oan211d1 U3083 ( .C1(n3828), .C2(n5187), .B(n5188), .A(n3958), .ZN(n5185) );
  oai222d1 U3084 ( .A1(n5190), .A2(n4431), .B1(n5191), .B2(n4431), .C1(n3821), 
        .C2(n5193), .ZN(n5183) );
  aoi21d1 U3085 ( .B1(n3823), .B2(n5195), .A(n5196), .ZN(n5191) );
  oai211d1 U3086 ( .C1(n5197), .C2(n5198), .A(n5199), .B(n5200), .ZN(n5195) );
  aoi31d1 U3087 ( .B1(n5201), .B2(n5202), .B3(n3830), .A(n3829), .ZN(n5200) );
  oai211d1 U3088 ( .C1(n3839), .C2(n5206), .A(n4698), .B(n5207), .ZN(n5202) );
  oai31d1 U3089 ( .B1(n5208), .B2(n5209), .B3(n5210), .A(n5211), .ZN(n5207) );
  oai222d1 U3090 ( .A1(n5212), .A2(n4409), .B1(n5665), .B2(n5214), .C1(
        images_bus[205]), .C2(n5215), .ZN(n5208) );
  oan211d1 U3092 ( .C1(n5217), .C2(n5218), .B(n5219), .A(n3897), .ZN(n5212) );
  aoi31d1 U3093 ( .B1(n3849), .B2(n5222), .B3(n5223), .A(n3846), .ZN(n5217) );
  aoim31d1 U3094 ( .B1(n5225), .B2(n5226), .B3(n5227), .A(n5228), .ZN(n5223)
         );
  aoi31d1 U3095 ( .B1(n5226), .B2(images_bus[209]), .B3(n5229), .A(n5230), 
        .ZN(n5228) );
  aoi321d1 U3096 ( .C1(n3875), .C2(n5232), .C3(n5233), .B1(n3875), .B2(n5234), 
        .A(n3852), .ZN(n5229) );
  aoi311d1 U3098 ( .C1(n5226), .C2(n5550), .C3(n5238), .A(n5239), .B(n5068), 
        .ZN(n5233) );
  aoi311d1 U3099 ( .C1(n5240), .C2(n5241), .C3(n3853), .A(n5068), .B(n5243), 
        .ZN(n5238) );
  oan211d1 U3100 ( .C1(images_bus[213]), .C2(n5244), .B(n5245), .A(n5246), 
        .ZN(n5243) );
  oai211d1 U3101 ( .C1(n5247), .C2(n5248), .A(n4315), .B(n5245), .ZN(n5241) );
  oan211d1 U3102 ( .C1(n5250), .C2(n5251), .B(n3869), .A(n5839), .ZN(n5247) );
  aoi31d1 U3103 ( .B1(n5253), .B2(n3896), .B3(n5255), .A(n5256), .ZN(n5250) );
  aoi31d1 U3104 ( .B1(n5257), .B2(n5258), .B3(n3857), .A(n5260), .ZN(n5255) );
  oai211d1 U3106 ( .C1(n5263), .C2(n5264), .A(n4954), .B(n5261), .ZN(n5258) );
  aoi31d1 U3107 ( .B1(n3810), .B2(n5267), .B3(n3721), .A(n3619), .ZN(n5263) );
  oai211d1 U3108 ( .C1(n5269), .C2(n5270), .A(n5271), .B(n5261), .ZN(n5267) );
  oan211d1 U3109 ( .C1(n5272), .C2(n5273), .B(n3734), .A(n5275), .ZN(n5269) );
  aoi311d1 U3110 ( .C1(n3699), .C2(n5277), .C3(n5748), .A(n5279), .B(n5280), 
        .ZN(n5272) );
  aon211d1 U3111 ( .C1(n3740), .C2(n5282), .B(n5283), .A(n3744), .ZN(n5277) );
  oan211d1 U3112 ( .C1(n5285), .C2(n5286), .B(images_bus[227]), .A(n5287), 
        .ZN(n5283) );
  oai211d1 U3113 ( .C1(n5288), .C2(n5289), .A(n5285), .B(n5290), .ZN(n5282) );
  oan211d1 U3114 ( .C1(n5291), .C2(n5292), .B(n3757), .A(n5294), .ZN(n5288) );
  aoim31d1 U3115 ( .B1(n5294), .B2(n5295), .B3(n5296), .A(n5297), .ZN(n5291)
         );
  aoim31d1 U3116 ( .B1(n3700), .B2(n5299), .B3(n5300), .A(n5301), .ZN(n5295)
         );
  aoi31d1 U3117 ( .B1(n5302), .B2(n5303), .B3(n5304), .A(n5305), .ZN(n5299) );
  aon211d1 U3118 ( .C1(n3801), .C2(n5307), .B(n5308), .A(n5309), .ZN(n5302) );
  aoi22d1 U3120 ( .A1(n5313), .A2(n3772), .B1(n3774), .B2(n5316), .ZN(n5311)
         );
  oan211d1 U3122 ( .C1(n5318), .C2(n5319), .B(n5544), .A(n5321), .ZN(n5313) );
  aoi211d1 U3123 ( .C1(n3777), .C2(n5323), .A(n5063), .B(n5324), .ZN(n5318) );
  oan211d1 U3124 ( .C1(n5325), .C2(n5326), .B(n5327), .A(n5328), .ZN(n5324) );
  oan211d1 U3125 ( .C1(n5329), .C2(n5330), .B(n5331), .A(n5332), .ZN(n5325) );
  aoi31d1 U3126 ( .B1(n5327), .B2(images_bus[249]), .B3(n5333), .A(n5334), 
        .ZN(n5329) );
  oan211d1 U3127 ( .C1(n5335), .C2(n5336), .B(n5337), .A(n5330), .ZN(n5333) );
  oai22d1 U3128 ( .A1(n5338), .A2(n5339), .B1(n5340), .B2(n4410), .ZN(n5336)
         );
  aoi211d1 U3129 ( .C1(n3788), .C2(n3577), .A(n5342), .B(n5343), .ZN(n5340) );
  aoi31d1 U3130 ( .B1(n3708), .B2(n5345), .B3(n5346), .A(n5347), .ZN(n5343) );
  aoi211d1 U3131 ( .C1(n5348), .C2(n5349), .A(n5350), .B(n5351), .ZN(n5346) );
  aon211d1 U3133 ( .C1(n3511), .C2(n3538), .B(n5356), .A(images_bus[257]), 
        .ZN(n5353) );
  oai211d1 U3135 ( .C1(n5360), .C2(n5361), .A(images_bus[271]), .B(n5362), 
        .ZN(n5357) );
  oan211d1 U3136 ( .C1(n5363), .C2(n3512), .B(n5365), .A(n5366), .ZN(n5361) );
  aoi21d1 U3139 ( .B1(n5372), .B2(n5373), .A(n5374), .ZN(n5369) );
  oai211d1 U3140 ( .C1(n5375), .C2(n5376), .A(n5377), .B(n5378), .ZN(n5372) );
  oan211d1 U3142 ( .C1(n5738), .C2(n3479), .B(n5381), .A(n5382), .ZN(n5376) );
  nd13d1 U3143 ( .A1(n5383), .A2(n5384), .A3(n5385), .ZN(n5381) );
  oai22d1 U3144 ( .A1(n5386), .A2(n3479), .B1(n5387), .B2(n5388), .ZN(n5385)
         );
  oai322d1 U3146 ( .C1(n5393), .C2(n5394), .C3(n5395), .A1(n5396), .A2(n3481), 
        .B1(n5398), .B2(n5391), .ZN(n5390) );
  aoi31d1 U3147 ( .B1(images_bus[299]), .B2(images_bus[298]), .B3(n5399), .A(
        n5400), .ZN(n5394) );
  aoi31d1 U3149 ( .B1(n3456), .B2(n3458), .B3(n5407), .A(n5408), .ZN(n5401) );
  oan211d1 U3150 ( .C1(n5409), .C2(n3453), .B(n5411), .A(n5412), .ZN(n5407) );
  aoi31d1 U3152 ( .B1(n3443), .B2(n5415), .B3(n5416), .A(n5417), .ZN(n5409) );
  oai31d1 U3153 ( .B1(n5418), .B2(n5419), .B3(n5420), .A(n5421), .ZN(n5415) );
  aoi311d1 U3154 ( .C1(n5422), .C2(n5423), .C3(n5424), .A(n5425), .B(n3480), 
        .ZN(n5419) );
  oai21d1 U3157 ( .B1(n5428), .B2(n5429), .A(n5430), .ZN(n5423) );
  aoi311d1 U3158 ( .C1(n3366), .C2(n5432), .C3(n3367), .A(n3337), .B(n3338), 
        .ZN(n5428) );
  aon211d1 U3159 ( .C1(n5436), .C2(n5437), .B(n5438), .A(n5439), .ZN(n5432) );
  oai211d1 U3161 ( .C1(n5444), .C2(n5445), .A(n5446), .B(n3335), .ZN(n5443) );
  oan211d1 U3163 ( .C1(n3336), .C2(n5450), .B(n5451), .A(n5452), .ZN(n5444) );
  aoi211d1 U3164 ( .C1(n5453), .C2(n5454), .A(n5455), .B(n3382), .ZN(n5450) );
  aon211d1 U3165 ( .C1(n5457), .C2(n3394), .B(n3336), .A(n3398), .ZN(n5453) );
  aoi21d1 U3166 ( .B1(n5460), .B2(n5461), .A(n5462), .ZN(n5457) );
  oan211d1 U3169 ( .C1(n5468), .C2(n5469), .B(n3271), .A(n5471), .ZN(n5467) );
  aoi211d1 U3170 ( .C1(n5472), .C2(n5473), .A(n5474), .B(n5475), .ZN(n5468) );
  aor211d1 U3171 ( .C1(n5476), .C2(n5472), .A(n5477), .B(n5478), .Z(n5473) );
  aon211d1 U3172 ( .C1(n5479), .C2(n5480), .B(n5481), .A(n3316), .ZN(n5476) );
  aoi21d1 U3173 ( .B1(n5483), .B2(n3253), .A(n5485), .ZN(n5479) );
  oai311d1 U3176 ( .C1(n5490), .C2(n5491), .C3(n5492), .A(n5493), .B(n5488), 
        .ZN(n5489) );
  aon211d1 U3177 ( .C1(n3312), .C2(n2808), .B(n5496), .A(n5497), .ZN(n5490) );
  oai211d1 U3178 ( .C1(n5498), .C2(n4304), .A(n3312), .B(n5499), .ZN(n5497) );
  aoi21d1 U3179 ( .B1(images_bus[374]), .B2(n5500), .A(n5501), .ZN(n5498) );
  aoim31d1 U3181 ( .B1(n5502), .B2(n5503), .B3(n5504), .A(n5496), .ZN(n5499)
         );
  aoi311d1 U3182 ( .C1(n5505), .C2(n3297), .C3(n5507), .A(n5496), .B(n5508), 
        .ZN(n5503) );
  oan211d1 U3183 ( .C1(n5509), .C2(n5510), .B(n5511), .A(n5512), .ZN(n5507) );
  aoi31d1 U3185 ( .B1(n5515), .B2(n5516), .B3(n5517), .A(n4638), .ZN(n5514) );
  aoi22d1 U3186 ( .A1(n3171), .A2(n5519), .B1(n3172), .B2(n5521), .ZN(n5517)
         );
  oai321d1 U3187 ( .C1(n3242), .C2(n5522), .C3(n3183), .B1(n5524), .B2(n5525), 
        .A(n5526), .ZN(n5519) );
  aoi311d1 U3190 ( .C1(n5529), .C2(n5530), .C3(n3188), .A(n5532), .B(n5533), 
        .ZN(n5522) );
  aoi21d1 U3191 ( .B1(n5534), .B2(n3189), .A(n5536), .ZN(n5533) );
  oai21d1 U3192 ( .B1(n4964), .B2(n5534), .A(n5537), .ZN(n5532) );
  aoim21d1 U3193 ( .B1(n5538), .B2(n4667), .A(n5539), .ZN(n5534) );
  oai211d1 U3194 ( .C1(n3140), .C2(n5541), .A(n3201), .B(n5543), .ZN(n5530) );
  aoi21d1 U3195 ( .B1(n3202), .B2(n5545), .A(n5546), .ZN(n5543) );
  aoi31d1 U3196 ( .B1(n5547), .B2(n3212), .B3(n5549), .A(n3203), .ZN(n5546) );
  aoi311d1 U3198 ( .C1(n5551), .C2(n5552), .C3(n3231), .A(n5553), .B(n3230), 
        .ZN(n5549) );
  oaim21d1 U3199 ( .B1(n5551), .B2(n5554), .A(n5555), .ZN(n5553) );
  aon211d1 U3200 ( .C1(n5556), .C2(n5551), .B(n5557), .A(n3223), .ZN(n5555) );
  aoi22d1 U3202 ( .A1(n3215), .A2(n5560), .B1(n5561), .B2(n5562), .ZN(n5547)
         );
  oai222d1 U3203 ( .A1(n5563), .A2(n4704), .B1(n5564), .B2(n5565), .C1(n5566), 
        .C2(n3027), .ZN(n5560) );
  oan211d1 U3204 ( .C1(n5568), .C2(n5569), .B(n3040), .A(n5571), .ZN(n5564) );
  aoim21d1 U3205 ( .B1(n4713), .B2(n4710), .A(n5572), .ZN(n5571) );
  oai22d1 U3207 ( .A1(n3026), .A2(n4720), .B1(n5574), .B2(n3046), .ZN(n5569)
         );
  aoi211d1 U3208 ( .C1(n4729), .C2(n5576), .A(n5577), .B(n4952), .ZN(n5574) );
  oai222d1 U3209 ( .A1(n5578), .A2(n3055), .B1(n5580), .B2(n3057), .C1(n3059), 
        .C2(n5583), .ZN(n5577) );
  aoi211d1 U3211 ( .C1(n3064), .C2(n5586), .A(n5587), .B(n5588), .ZN(n5580) );
  aoi21d1 U3212 ( .B1(n3065), .B2(n5589), .A(n5590), .ZN(n5588) );
  oai211d1 U3213 ( .C1(n3073), .C2(n5592), .A(n5593), .B(n5594), .ZN(n5586) );
  aoi221d1 U3215 ( .B1(n5599), .B2(n3117), .C1(n5596), .C2(n5600), .A(n5601), 
        .ZN(n5598) );
  oai221d1 U3216 ( .B1(n5602), .B2(n5603), .C1(n3082), .C2(n5605), .A(n5606), 
        .ZN(n5601) );
  ora211d1 U3217 ( .C1(n4301), .C2(n3087), .A(n5608), .B(n5609), .Z(n5605) );
  oan211d1 U3218 ( .C1(n4757), .C2(n5610), .B(n5611), .A(n5612), .ZN(n5609) );
  oan211d1 U3219 ( .C1(n5613), .C2(n5614), .B(n5615), .A(n5616), .ZN(n5612) );
  aoi22d1 U3220 ( .A1(n3015), .A2(n5618), .B1(n5619), .B2(n5620), .ZN(n5615)
         );
  oai211d1 U3221 ( .C1(n2929), .C2(n4785), .A(n5622), .B(n5623), .ZN(n5618) );
  aoi311d1 U3222 ( .C1(n5624), .C2(n4788), .C3(n2925), .A(n2923), .B(n5627), 
        .ZN(n5623) );
  oan211d1 U3224 ( .C1(n5629), .C2(n5630), .B(n2924), .A(n5632), .ZN(n5622) );
  aoi21d1 U3225 ( .B1(n5613), .B2(n2935), .A(n2926), .ZN(n5632) );
  oai21d1 U3227 ( .B1(n3007), .B2(n2929), .A(n5637), .ZN(n5630) );
  oai22d1 U3228 ( .A1(n5638), .A2(n5639), .B1(n5640), .B2(n5641), .ZN(n5629)
         );
  aoim211d1 U3229 ( .C1(n5638), .C2(n2955), .A(n5643), .B(n2952), .ZN(n5640)
         );
  oai22d1 U3230 ( .A1(n5645), .A2(n4807), .B1(n5646), .B2(n2954), .ZN(n5643)
         );
  aoi211d1 U3231 ( .C1(n2991), .C2(n5649), .A(n5650), .B(n5651), .ZN(n5645) );
  oai22d1 U3232 ( .A1(n5646), .A2(n2997), .B1(n5653), .B2(n5654), .ZN(n5650)
         );
  aoi211d1 U3233 ( .C1(n2961), .C2(n5649), .A(n5656), .B(n5657), .ZN(n5653) );
  oai22d1 U3234 ( .A1(n5658), .A2(n5659), .B1(n5660), .B2(n5661), .ZN(n5656)
         );
  aoi211d1 U3235 ( .C1(n5662), .C2(n5663), .A(n5664), .B(n2972), .ZN(n5660) );
  oai22d1 U3236 ( .A1(n5658), .A2(n5666), .B1(n5667), .B2(n5668), .ZN(n5664)
         );
  aoi221d1 U3237 ( .B1(n2978), .B2(n5670), .C1(n5671), .C2(n5663), .A(n5672), 
        .ZN(n5667) );
  oai22d1 U3238 ( .A1(n5673), .A2(n4929), .B1(n5674), .B2(n5675), .ZN(n5670)
         );
  aoi321d1 U3239 ( .C1(n2851), .C2(n5677), .C3(n5678), .B1(n5679), .B2(n5680), 
        .A(n5681), .ZN(n5673) );
  oai21d1 U3240 ( .B1(n4930), .B2(n5674), .A(n5682), .ZN(n5681) );
  oai211d1 U3241 ( .C1(n2838), .C2(n4870), .A(n2853), .B(n5685), .ZN(n5680) );
  aoi22d1 U3242 ( .A1(n2855), .A2(n5686), .B1(n2856), .B2(n5688), .ZN(n5685)
         );
  oai211d1 U3243 ( .C1(n2837), .C2(n2870), .A(n2867), .B(n5692), .ZN(n5688) );
  aoi22d1 U3244 ( .A1(n2869), .A2(n5694), .B1(n4878), .B2(n5695), .ZN(n5692)
         );
  oaim211d1 U3245 ( .C1(n5695), .C2(n4879), .A(n4885), .B(n5696), .ZN(n5694)
         );
  aon211d1 U3269 ( .C1(n5572), .C2(n5729), .B(n4721), .A(n3048), .ZN(n5568) );
  aoim211d1 U3271 ( .C1(n4702), .C2(n5566), .A(n5707), .B(n4705), .ZN(n5563)
         );
  nd13d1 U3308 ( .A1(n4483), .A2(n5735), .A3(n5375), .ZN(n5391) );
  aoi31d1 U3337 ( .B1(n3881), .B2(n5760), .B3(n3880), .A(n5764), .ZN(n5197) );
  aoi22d1 U3343 ( .A1(n5770), .A2(n7243), .B1(n3826), .B2(n5749), .ZN(n5190)
         );
  oai21d1 U3346 ( .B1(n5774), .B2(n5169), .A(n3945), .ZN(n5174) );
  aoi211d1 U3363 ( .C1(n5787), .C2(images_bus[64]), .A(n5008), .B(n5021), .ZN(
        N26364) );
  aoi22d1 U3368 ( .A1(n4196), .A2(n5801), .B1(n4199), .B2(n5803), .ZN(n5787)
         );
  oai21d1 U3369 ( .B1(n5804), .B2(n5805), .A(n5778), .ZN(n5801) );
  oai22d1 U3371 ( .A1(images_bus[69]), .A2(n5810), .B1(n5811), .B2(n5812), 
        .ZN(n5808) );
  oan211d1 U3372 ( .C1(n5813), .C2(n5814), .B(n5033), .A(n6641), .ZN(n5811) );
  or03d0 U3373 ( .A1(n5815), .A2(n6641), .A3(n5298), .Z(n5814) );
  oai211d1 U3374 ( .C1(images_bus[71]), .C2(n5816), .A(n5817), .B(n5778), .ZN(
        n5813) );
  aon211d1 U3375 ( .C1(n4182), .C2(n5819), .B(n5820), .A(n5821), .ZN(n5817) );
  oai211d1 U3376 ( .C1(n5822), .C2(n5823), .A(n5824), .B(n4747), .ZN(n5819) );
  aon211d1 U3377 ( .C1(n4152), .C2(n5827), .B(n5691), .A(n5828), .ZN(n5824) );
  aoi211d1 U3378 ( .C1(n5829), .C2(n5830), .A(n5204), .B(n5827), .ZN(n5822) );
  oai211d1 U3379 ( .C1(n5831), .C2(n5832), .A(n4156), .B(n4746), .ZN(n5830) );
  aon211d1 U3380 ( .C1(n4157), .C2(n5836), .B(n4503), .A(n4180), .ZN(n5832) );
  oai211d1 U3381 ( .C1(n5838), .C2(n4177), .A(n4746), .B(n5840), .ZN(n5836) );
  oan211d1 U3384 ( .C1(n5845), .C2(n4174), .B(n5847), .A(n5848), .ZN(n5843) );
  aoi211d1 U3385 ( .C1(n4175), .C2(n5106), .A(n5850), .B(n4506), .ZN(n5845) );
  oai22d1 U3387 ( .A1(n5852), .A2(n5853), .B1(n5854), .B2(n4158), .ZN(n5850)
         );
  oan211d1 U3388 ( .C1(n5856), .C2(n5857), .B(n4163), .A(n4326), .ZN(n5854) );
  oai22d1 U3389 ( .A1(images_bus[87]), .A2(n5859), .B1(n5860), .B2(n5861), 
        .ZN(n5857) );
  aoi31d1 U3390 ( .B1(n4169), .B2(n5863), .B3(N9106), .A(n4324), .ZN(n5860) );
  oai211d1 U3392 ( .C1(n5865), .C2(n5866), .A(n5867), .B(n5868), .ZN(n5863) );
  aon211d1 U3393 ( .C1(n5869), .C2(n4170), .B(n5871), .A(n5872), .ZN(n5867) );
  oan211d1 U3394 ( .C1(n5873), .C2(n5874), .B(n5875), .A(n5876), .ZN(n5869) );
  oai222d1 U3396 ( .A1(n5880), .A2(n5881), .B1(n5882), .B2(n5883), .C1(n5884), 
        .C2(n5885), .ZN(n5877) );
  aon211d1 U3397 ( .C1(n5886), .C2(n5887), .B(n6948), .A(n5888), .ZN(n5883) );
  oai211d1 U3399 ( .C1(n5892), .C2(n5893), .A(n4066), .B(n5895), .ZN(n5891) );
  oan211d1 U3400 ( .C1(n5896), .C2(n5897), .B(n4124), .A(n5899), .ZN(n5892) );
  oan211d1 U3401 ( .C1(n5900), .C2(n5901), .B(n4071), .A(n6056), .ZN(n5896) );
  aoi31d1 U3402 ( .B1(images_bus[105]), .B2(n5903), .B3(n4123), .A(n5905), 
        .ZN(n5900) );
  aon211d1 U3403 ( .C1(n4075), .C2(n5907), .B(n5908), .A(n5909), .ZN(n5903) );
  oai21d1 U3405 ( .B1(n6576), .B2(n5913), .A(n5914), .ZN(n5912) );
  oai22d1 U3406 ( .A1(images_bus[109]), .A2(n5915), .B1(n5916), .B2(n5917), 
        .ZN(n5913) );
  oai22d1 U3409 ( .A1(n5922), .A2(n5923), .B1(n5924), .B2(n5026), .ZN(n5919)
         );
  oan211d1 U3410 ( .C1(n5925), .C2(n5926), .B(n4082), .A(n5575), .ZN(n5924) );
  aoi31d1 U3411 ( .B1(images_bus[115]), .B2(n5928), .B3(n5929), .A(n5930), 
        .ZN(n5925) );
  oai211d1 U3412 ( .C1(n4101), .C2(n5932), .A(n4102), .B(N9484), .ZN(n5928) );
  aon211d1 U3413 ( .C1(images_bus[117]), .C2(n5934), .B(n5935), .A(n5929), 
        .ZN(n5932) );
  oai31d1 U3414 ( .B1(n5936), .B2(n4090), .B3(n5938), .A(n4087), .ZN(n5934) );
  aoi31d1 U3416 ( .B1(n5941), .B2(n5942), .B3(n5943), .A(n5030), .ZN(n5938) );
  aon211d1 U3417 ( .C1(n4095), .C2(n5945), .B(n5946), .A(n5024), .ZN(n5942) );
  oai321d1 U3418 ( .C1(n5947), .C2(n5948), .C3(n3998), .B1(n5950), .B2(n5951), 
        .A(n3984), .ZN(n5945) );
  oai21d1 U3420 ( .B1(n5041), .B2(images_bus[127]), .A(n5954), .ZN(n5953) );
  aon211d1 U3421 ( .C1(n5955), .C2(N9696), .B(n5956), .A(n4003), .ZN(n5947) );
  oan211d1 U3422 ( .C1(n3997), .C2(n4009), .B(n5960), .A(n5961), .ZN(n5955) );
  aon211d1 U3423 ( .C1(n5962), .C2(n4015), .B(n5963), .A(n4012), .ZN(n5960) );
  aoi221d1 U3428 ( .B1(n5969), .B2(n5970), .C1(n5971), .C2(n5081), .A(n5972), 
        .ZN(n5966) );
  oai211d1 U3430 ( .C1(n5977), .C2(n5978), .A(n4045), .B(n4029), .ZN(n5974) );
  oan211d1 U3431 ( .C1(n5981), .C2(n3974), .B(n5983), .A(n5984), .ZN(n5978) );
  oai211d1 U3432 ( .C1(n5985), .C2(n5986), .A(n3966), .B(n3911), .ZN(n5983) );
  oan211d1 U3433 ( .C1(n5144), .C2(n5989), .B(n5990), .A(n4424), .ZN(n5986) );
  oai21d1 U3436 ( .B1(n5995), .B2(n5989), .A(n5996), .ZN(n5991) );
  oai22d1 U3438 ( .A1(n5999), .A2(n6000), .B1(n6001), .B2(n6002), .ZN(n5998)
         );
  aon211d1 U3440 ( .C1(n3951), .C2(n6005), .B(n6006), .A(n3953), .ZN(n6001) );
  oai22d1 U3442 ( .A1(n5193), .A2(n6008), .B1(n6009), .B2(n6010), .ZN(n6005)
         );
  aon211d1 U3443 ( .C1(n5770), .C2(n6011), .B(n6012), .A(n3821), .ZN(n6010) );
  oan211d1 U3444 ( .C1(n6013), .C2(n6014), .B(n6015), .A(n6016), .ZN(n6012) );
  oai31d1 U3445 ( .B1(n6011), .B2(n6017), .B3(n5749), .A(n3824), .ZN(n6015) );
  aoi31d1 U3447 ( .B1(n6019), .B2(n6020), .B3(n6021), .A(n6022), .ZN(n6017) );
  oan211d1 U3448 ( .C1(n6023), .C2(n3898), .B(n3831), .A(n6934), .ZN(n6021) );
  aoi221d1 U3451 ( .B1(n6031), .B2(n6032), .C1(n3836), .C2(n6034), .A(n6035), 
        .ZN(n6027) );
  oai211d1 U3452 ( .C1(n6036), .C2(n5214), .A(n6037), .B(n3842), .ZN(n6032) );
  aor31d1 U3454 ( .B1(n2800), .B2(n6036), .B3(n6040), .A(n4409), .Z(n6037) );
  oai22d1 U3456 ( .A1(n6042), .A2(n6043), .B1(n6044), .B2(n3848), .ZN(n6041)
         );
  aoi22d1 U3457 ( .A1(n6046), .A2(n6047), .B1(n3853), .B2(n6048), .ZN(n6042)
         );
  oai211d1 U3458 ( .C1(n6049), .C2(n6050), .A(n3899), .B(n6052), .ZN(n6048) );
  aoi221d1 U3459 ( .B1(n6053), .B2(n6054), .C1(n6055), .C2(n3618), .A(n6057), 
        .ZN(n6049) );
  oai22d1 U3460 ( .A1(n6058), .A2(n6059), .B1(n6060), .B2(n3723), .ZN(n6054)
         );
  aoi22d1 U3462 ( .A1(n6063), .A2(n6064), .B1(n3734), .B2(n6065), .ZN(n6060)
         );
  aon211d1 U3464 ( .C1(images_bus[227]), .C2(n6067), .B(n5287), .A(n6068), 
        .ZN(n6064) );
  aor31d1 U3465 ( .B1(n6068), .B2(n6069), .B3(n5274), .A(n5286), .Z(n6067) );
  aon211d1 U3466 ( .C1(n6071), .C2(n3748), .B(n4691), .A(n6073), .ZN(n6069) );
  aor311d1 U3467 ( .C1(n3759), .C2(n3757), .C3(n6075), .A(n6076), .B(n6077), 
        .Z(n6071) );
  aoi31d1 U3468 ( .B1(n6078), .B2(n5655), .B3(n6080), .A(n6081), .ZN(n6075) );
  aoi21d1 U3469 ( .B1(n6082), .B2(n3764), .A(n3679), .ZN(n6081) );
  oan211d1 U3471 ( .C1(n6085), .C2(n5173), .B(n3805), .A(n5648), .ZN(n6080) );
  aoi31d1 U3473 ( .B1(n6078), .B2(n6086), .B3(n6087), .A(n6088), .ZN(n6085) );
  aon211d1 U3474 ( .C1(n3802), .C2(n6090), .B(n6091), .A(n5309), .ZN(n6086) );
  oai22d1 U3475 ( .A1(images_bus[239]), .A2(n6092), .B1(n6093), .B2(n6094), 
        .ZN(n6090) );
  oan211d1 U3476 ( .C1(n6095), .C2(n6096), .B(n3800), .A(n3692), .ZN(n6093) );
  aon211d1 U3477 ( .C1(n6099), .C2(n3779), .B(n6101), .A(n6102), .ZN(n6096) );
  aoi211d1 U3478 ( .C1(n6103), .C2(n6104), .A(n6105), .B(n6106), .ZN(n6101) );
  aon211d1 U3479 ( .C1(n6107), .C2(n6108), .B(n6109), .A(n6110), .ZN(n6104) );
  aoi21d1 U3480 ( .B1(n6111), .B2(n6112), .A(n3681), .ZN(n6107) );
  aon211d1 U3483 ( .C1(n3521), .C2(n6118), .B(n3573), .A(n6120), .ZN(n6116) );
  oai211d1 U3484 ( .C1(n6121), .C2(n6122), .A(images_bus[253]), .B(n3684), 
        .ZN(n6120) );
  aoi211d1 U3485 ( .C1(n5348), .C2(n6124), .A(n6125), .B(n6126), .ZN(n6121) );
  oan211d1 U3486 ( .C1(n6127), .C2(n6128), .B(n6129), .A(n6130), .ZN(n6126) );
  aoi22d1 U3487 ( .A1(n6131), .A2(n6132), .B1(n3520), .B2(n6134), .ZN(n6127)
         );
  aoi211d1 U3488 ( .C1(n6135), .C2(n6136), .A(n6137), .B(n3564), .ZN(n6132) );
  oan211d1 U3490 ( .C1(n6142), .C2(n6143), .B(n6144), .A(n6145), .ZN(n6141) );
  oai321d1 U3493 ( .C1(n6150), .C2(n7016), .C3(n5410), .B1(n6151), .B2(n3518), 
        .A(n6153), .ZN(n6149) );
  oan211d1 U3495 ( .C1(n6158), .C2(n3518), .B(n6159), .A(n12149), .ZN(n6156)
         );
  aoi21d1 U3497 ( .B1(n6163), .B2(n6164), .A(n6165), .ZN(n6161) );
  oan211d1 U3499 ( .C1(n6169), .C2(n3504), .B(n6171), .A(n6172), .ZN(n6168) );
  oan211d1 U3501 ( .C1(n5404), .C2(n6177), .B(n6178), .A(n6169), .ZN(n6175) );
  oan211d1 U3503 ( .C1(n6181), .C2(n6177), .B(n6182), .A(n6183), .ZN(n6180) );
  oai31d1 U3505 ( .B1(n6187), .B2(n6188), .B3(n3442), .A(n6190), .ZN(n6186) );
  oai211d1 U3506 ( .C1(n6191), .C2(n6192), .A(n6193), .B(n6194), .ZN(n6187) );
  aoi211d1 U3507 ( .C1(n6195), .C2(n6196), .A(n6197), .B(n6198), .ZN(n6192) );
  aoi22d1 U3508 ( .A1(n3419), .A2(n5737), .B1(n3365), .B2(n6201), .ZN(n6195)
         );
  oai211d1 U3509 ( .C1(n6202), .C2(n6203), .A(n6204), .B(n6205), .ZN(n6201) );
  aoi211d1 U3510 ( .C1(n6206), .C2(n3413), .A(n6208), .B(n3415), .ZN(n6202) );
  aoi31d1 U3512 ( .B1(n4668), .B2(n6211), .B3(n3356), .A(n6213), .ZN(n6206) );
  oai321d1 U3515 ( .C1(n6214), .C2(n6217), .C3(n4989), .B1(n3373), .B2(n6004), 
        .A(n3411), .ZN(n6211) );
  oai21d1 U3516 ( .B1(n6216), .B2(n6219), .A(n6220), .ZN(n6214) );
  oai31d1 U3517 ( .B1(n6221), .B2(n6222), .B3(n6223), .A(n6224), .ZN(n6219) );
  aon211d1 U3518 ( .C1(n5634), .C2(n5445), .B(n6226), .A(n6227), .ZN(n6224) );
  oai211d1 U3519 ( .C1(n6228), .C2(n3400), .A(n6230), .B(n6231), .ZN(n6221) );
  aoi211d1 U3520 ( .C1(n6232), .C2(n5927), .A(n6233), .B(n6234), .ZN(n6228) );
  aoi31d1 U3521 ( .B1(n3359), .B2(n5724), .B3(n6236), .A(n6237), .ZN(n6234) );
  oan211d1 U3522 ( .C1(n6238), .C2(n6239), .B(n3377), .A(n6241), .ZN(n6236) );
  aoi31d1 U3523 ( .B1(n3358), .B2(n6243), .B3(n6244), .A(n6245), .ZN(n6238) );
  aoi31d1 U3524 ( .B1(n3383), .B2(n6247), .B3(n6248), .A(n6249), .ZN(n6245) );
  aoi31d1 U3525 ( .B1(n2801), .B2(n3398), .B3(n6251), .A(n6252), .ZN(n6248) );
  aoim211d1 U3526 ( .C1(n6253), .C2(n2801), .A(n6254), .B(n6249), .ZN(n6244)
         );
  aon211d1 U3529 ( .C1(n6256), .C2(n6257), .B(n6258), .A(images_bus[341]), 
        .ZN(n6255) );
  aoi21d1 U3530 ( .B1(n3397), .B2(n5825), .A(n6260), .ZN(n6256) );
  aoi31d1 U3531 ( .B1(n6257), .B2(n5721), .B3(n6261), .A(n6262), .ZN(n6260) );
  aoi22d1 U3532 ( .A1(n6263), .A2(n5397), .B1(n3387), .B2(n6265), .ZN(n6261)
         );
  oai211d1 U3533 ( .C1(n6266), .C2(n3391), .A(n3392), .B(n6269), .ZN(n6265) );
  aoi321d1 U3534 ( .C1(n3270), .C2(n6271), .C3(n6272), .B1(n3389), .B2(n3268), 
        .A(n6274), .ZN(n6266) );
  aoi31d1 U3536 ( .B1(n3357), .B2(n6277), .B3(n6278), .A(n6275), .ZN(n6272) );
  aoi321d1 U3537 ( .C1(n3272), .C2(n6280), .C3(n3273), .B1(n3272), .B2(n6097), 
        .A(n6281), .ZN(n6278) );
  aon211d1 U3538 ( .C1(images_bus[352]), .C2(n5475), .B(n6282), .A(n6283), 
        .ZN(n6280) );
  oai21d1 U3540 ( .B1(n5252), .B2(n4586), .A(n3327), .ZN(n6285) );
  aoi31d1 U3541 ( .B1(n6288), .B2(n6289), .B3(n6290), .A(n3324), .ZN(n6284) );
  aoi211d1 U3543 ( .C1(n3318), .C2(n5988), .A(n6286), .B(n6294), .ZN(n6290) );
  aoi21d1 U3544 ( .B1(n6295), .B2(n6296), .A(n3276), .ZN(n6289) );
  aon211d1 U3547 ( .C1(n4977), .C2(n3314), .B(n6304), .A(n3315), .ZN(n6300) );
  oai21d1 U3549 ( .B1(n6307), .B2(n6308), .A(n6309), .ZN(n6304) );
  aon211d1 U3551 ( .C1(n6311), .C2(n6312), .B(n6313), .A(n6314), .ZN(n6308) );
  oai31d1 U3552 ( .B1(n6315), .B2(n4610), .B3(n6307), .A(n6316), .ZN(n6312) );
  or02d0 U3553 ( .A1(n6317), .A2(n6318), .Z(n4610) );
  oai21d1 U3554 ( .B1(n6319), .B2(n6320), .A(n6321), .ZN(n6315) );
  oai321d1 U3555 ( .C1(n6322), .C2(n5491), .C3(n6323), .B1(n3291), .B2(n5523), 
        .A(n5487), .ZN(n6321) );
  aon211d1 U3556 ( .C1(n6325), .C2(n6326), .B(n5492), .A(n6327), .ZN(n6322) );
  oai21d1 U3557 ( .B1(n3308), .B2(n5716), .A(n6329), .ZN(n6325) );
  aon211d1 U3558 ( .C1(n2802), .C2(n6331), .B(n6332), .A(n3308), .ZN(n6329) );
  aoi21d1 U3559 ( .B1(n6333), .B2(n6334), .A(n6335), .ZN(n6332) );
  oai21d1 U3561 ( .B1(images_bus[375]), .B2(n5500), .A(n6336), .ZN(n6334) );
  oai211d1 U3562 ( .C1(n6337), .C2(n6338), .A(n6331), .B(n6339), .ZN(n6336) );
  aoi31d1 U3563 ( .B1(n6340), .B2(n6341), .B3(n6342), .A(n6343), .ZN(n6339) );
  oan211d1 U3564 ( .C1(n3301), .C2(n5370), .B(n3302), .A(n6346), .ZN(n6343) );
  aon211d1 U3565 ( .C1(images_bus[379]), .C2(n6341), .B(n6347), .A(n3300), 
        .ZN(n6338) );
  oai31d1 U3566 ( .B1(n6337), .B2(n6349), .B3(n4902), .A(n6340), .ZN(n6341) );
  aoi311d1 U3567 ( .C1(n6350), .C2(n6351), .C3(n6352), .A(n6353), .B(n6354), 
        .ZN(n6349) );
  oan211d1 U3568 ( .C1(n3168), .C2(n3138), .B(n3297), .A(n3254), .ZN(n6354) );
  aoi321d1 U3570 ( .C1(n6357), .C2(n3163), .C3(n6359), .B1(n3167), .B2(n6361), 
        .A(n6362), .ZN(n6352) );
  oan211d1 U3573 ( .C1(n3141), .C2(n6367), .B(n7604), .A(n6369), .ZN(n6357) );
  aoim31d1 U3574 ( .B1(n6370), .B2(n3245), .B3(n6372), .A(n6361), .ZN(n6369)
         );
  aoi31d1 U3575 ( .B1(n3243), .B2(n6373), .B3(n6374), .A(n6361), .ZN(n6370) );
  aoi311d1 U3576 ( .C1(n6375), .C2(n6376), .C3(n6373), .A(n6377), .B(n6378), 
        .ZN(n6374) );
  or03d0 U3577 ( .A1(n6379), .A2(n6380), .A3(n6381), .Z(n6375) );
  aon211d1 U3578 ( .C1(n6382), .C2(n3186), .B(n6384), .A(N13762), .ZN(n6381)
         );
  aor22d1 U3579 ( .A1(n6385), .A2(n6386), .B1(n6387), .B2(n3142), .Z(n6382) );
  oan211d1 U3580 ( .C1(n3193), .C2(n5906), .B(n3241), .A(n6391), .ZN(n6387) );
  aoi21d1 U3581 ( .B1(n6392), .B2(n6393), .A(n6394), .ZN(n6385) );
  oai22d1 U3584 ( .A1(n3205), .A2(n5506), .B1(n6401), .B2(n6402), .ZN(n6396)
         );
  oai31d1 U3586 ( .B1(n6405), .B2(n6406), .B3(n6407), .A(n6408), .ZN(n6404) );
  oai211d1 U3587 ( .C1(n6409), .C2(n6410), .A(n3238), .B(n6412), .ZN(n6408) );
  oai22d1 U3588 ( .A1(n3208), .A2(n4302), .B1(n6414), .B2(n6415), .ZN(n6410)
         );
  aoim31d1 U3589 ( .B1(n6416), .B2(N13986), .B3(n6417), .A(n6417), .ZN(n6414)
         );
  aon211d1 U3590 ( .C1(n6418), .C2(n6419), .B(n6420), .A(n3208), .ZN(n6405) );
  aon211d1 U3592 ( .C1(n3029), .C2(n6426), .B(n6427), .A(n3224), .ZN(n6422) );
  aon211d1 U3594 ( .C1(n6432), .C2(n6433), .B(n6434), .A(n6435), .ZN(n6426) );
  aoi31d1 U3595 ( .B1(n6436), .B2(n3130), .B3(n6438), .A(n6439), .ZN(n6435) );
  aoim21d1 U3596 ( .B1(n6440), .B2(n6441), .A(n6429), .ZN(n6439) );
  oan211d1 U3597 ( .C1(n12140), .C2(n6442), .B(n3051), .A(n6434), .ZN(n6438)
         );
  oai22d1 U3600 ( .A1(n6447), .A2(n6448), .B1(n6444), .B2(n6449), .ZN(n6446)
         );
  aon211d1 U3601 ( .C1(images_bus[421]), .C2(n4729), .B(n6448), .A(n6599), 
        .ZN(n6449) );
  aoi211d1 U3602 ( .C1(n6450), .C2(n6451), .A(n6452), .B(n6453), .ZN(n6447) );
  oai22d1 U3604 ( .A1(n6456), .A2(n6457), .B1(n6458), .B2(n6459), .ZN(n6452)
         );
  aoim31d1 U3605 ( .B1(n6460), .B2(N14322), .B3(n6457), .A(n6461), .ZN(n6458)
         );
  aoi211d1 U3606 ( .C1(n6462), .C2(n6463), .A(n6464), .B(n6465), .ZN(n6461) );
  oai322d1 U3608 ( .C1(n6468), .C2(n3078), .C3(n6470), .A1(n6471), .A2(n6472), 
        .B1(n6473), .B2(n6474), .ZN(n6467) );
  aoi22d1 U3609 ( .A1(n3094), .A2(n6476), .B1(n6477), .B2(n6478), .ZN(n6473)
         );
  oai222d1 U3610 ( .A1(n6479), .A2(n6480), .B1(n3131), .B2(n6482), .C1(n6483), 
        .C2(n3107), .ZN(n6476) );
  aon211d1 U3612 ( .C1(images_bus[439]), .C2(n6486), .B(n6487), .A(
        images_bus[438]), .ZN(n6482) );
  aoim31d1 U3614 ( .B1(n3101), .B2(n12167), .B3(n6483), .A(n6489), .ZN(n6479)
         );
  oan211d1 U3615 ( .C1(n6483), .C2(n6490), .B(n6491), .A(n6492), .ZN(n6489) );
  aon211d1 U3616 ( .C1(n6493), .C2(n6494), .B(n6495), .A(n3095), .ZN(n6491) );
  oan211d1 U3617 ( .C1(n6497), .C2(n4774), .B(n6498), .A(n6499), .ZN(n6495) );
  aoi211d1 U3620 ( .C1(n6503), .C2(n6504), .A(n6505), .B(n6506), .ZN(n6497) );
  oan211d1 U3621 ( .C1(n3011), .C2(n6083), .B(n2927), .A(n6509), .ZN(n6506) );
  aon211d1 U3622 ( .C1(n6510), .C2(n6511), .B(n5635), .A(n5628), .ZN(n6505) );
  oai211d1 U3624 ( .C1(n2955), .C2(n6514), .A(n6515), .B(n6516), .ZN(n6513) );
  aoi22d1 U3625 ( .A1(n6517), .A2(n6518), .B1(n2953), .B2(n6520), .ZN(n6516)
         );
  oai211d1 U3626 ( .C1(n6521), .C2(n6522), .A(n2965), .B(n6524), .ZN(n6520) );
  aoi22d1 U3627 ( .A1(n2989), .A2(n6526), .B1(n6527), .B2(n6518), .ZN(n6524)
         );
  oai211d1 U3628 ( .C1(n6521), .C2(n6528), .A(n2963), .B(n6530), .ZN(n6526) );
  aoi22d1 U3629 ( .A1(n2959), .A2(n6532), .B1(n2960), .B2(n6534), .ZN(n6530)
         );
  oaim211d1 U3631 ( .C1(n6535), .C2(n5662), .A(n6536), .B(n6537), .ZN(n6532)
         );
  aoi22d1 U3632 ( .A1(n2971), .A2(n6539), .B1(n6534), .B2(n2970), .ZN(n6537)
         );
  oai221d1 U3634 ( .B1(n6541), .B2(n6542), .C1(n2920), .C2(n4934), .A(n2818), 
        .ZN(n6539) );
  aoi211d1 U3636 ( .C1(n6535), .C2(n4850), .A(n6545), .B(n4852), .ZN(n6541) );
  oai21d1 U3637 ( .B1(n4929), .B2(n6546), .A(n2825), .ZN(n4852) );
  oai322d1 U3638 ( .C1(n4929), .C2(n2832), .C3(n6549), .A1(n2805), .A2(n4856), 
        .B1(n2832), .B2(n4857), .ZN(n6545) );
  aoi21d1 U3649 ( .B1(n4791), .B2(n6504), .A(n2942), .ZN(n6510) );
  oai21d1 U3650 ( .B1(n6083), .B2(n6509), .A(images_bus[448]), .ZN(n6504) );
  oan211d1 U3653 ( .C1(n3105), .C2(n6428), .B(n3102), .A(n6557), .ZN(n6493) );
  aon211d1 U3654 ( .C1(n5344), .C2(n6557), .B(n6559), .A(n3108), .ZN(n6490) );
  aon211d1 U3657 ( .C1(images_bus[435]), .C2(n6563), .B(n6564), .A(n3081), 
        .ZN(n6472) );
  oai21d1 U3660 ( .B1(n6569), .B2(n6570), .A(n3132), .ZN(n6462) );
  oai22d1 U3663 ( .A1(n3075), .A2(n4406), .B1(n3121), .B2(n6573), .ZN(n6570)
         );
  oan211d1 U3667 ( .C1(n3058), .C2(n5980), .B(n3054), .A(n4729), .ZN(n6450) );
  aon211d1 U3668 ( .C1(n5729), .C2(n6577), .B(n6578), .A(n6574), .ZN(n6432) );
  oai211d1 U3671 ( .C1(n6580), .C2(n6993), .A(n6581), .B(n6582), .ZN(n6419) );
  aoi31d1 U3672 ( .B1(n6583), .B2(n6584), .B3(n6585), .A(n3221), .ZN(n6582) );
  aoi31d1 U3674 ( .B1(n5364), .B2(n6587), .B3(n6583), .A(n6588), .ZN(n6580) );
  or03d0 U3685 ( .A1(n6595), .A2(n6346), .A3(n6335), .Z(n6337) );
  nd13d1 U3686 ( .A1(n6323), .A2(n4305), .A3(n5044), .ZN(n6335) );
  aoi21d1 U3706 ( .B1(images_bus[319]), .B2(n6191), .A(n7232), .ZN(n6196) );
  nd13d1 U3708 ( .A1(n6177), .A2(n4994), .A3(n5833), .ZN(n6190) );
  aon211d1 U3743 ( .C1(n3880), .C2(n6035), .B(n12170), .A(n3830), .ZN(n6019)
         );
  oai21d1 U3748 ( .B1(n6119), .B2(n6008), .A(images_bus[192]), .ZN(n6011) );
  aoi21d1 U3769 ( .B1(images_bus[127]), .B2(n5950), .A(n5053), .ZN(n5956) );
  aoim2m11d1 U3790 ( .C1(n6668), .C2(n6669), .B(n5795), .A(n5008), .ZN(N26363)
         );
  aoim21d1 U3795 ( .B1(n6684), .B2(n6685), .A(n6686), .ZN(n6669) );
  aoi31d1 U3796 ( .B1(n6687), .B2(n6688), .B3(n6689), .A(n6690), .ZN(n6684) );
  aoi22d1 U3797 ( .A1(n6691), .A2(n6692), .B1(n4239), .B2(n6694), .ZN(n6689)
         );
  oai211d1 U3798 ( .C1(n6695), .C2(n6696), .A(n6697), .B(n5306), .ZN(n6692) );
  aoi21d1 U3799 ( .B1(n4244), .B2(n6700), .A(n4246), .ZN(n6695) );
  oai31d1 U3801 ( .B1(n6704), .B2(n6705), .B3(n6706), .A(n4274), .ZN(n6703) );
  oai222d1 U3802 ( .A1(n6708), .A2(n5800), .B1(n6709), .B2(n6710), .C1(
        images_bus[42]), .C2(n6711), .ZN(n6704) );
  aoi211d1 U3806 ( .C1(n6721), .C2(n6722), .A(n4257), .B(n6724), .ZN(n6717) );
  oai21d1 U3807 ( .B1(n6725), .B2(n6726), .A(n6727), .ZN(n6716) );
  aon211d1 U3808 ( .C1(n6728), .C2(n6729), .B(n6730), .A(n4514), .ZN(n6726) );
  aoi221d1 U3809 ( .B1(n4264), .B2(n6733), .C1(n6734), .C2(n6735), .A(n4265), 
        .ZN(n6729) );
  aoi211d1 U3810 ( .C1(n4215), .C2(n6738), .A(n6739), .B(n6740), .ZN(n6728) );
  oai211d1 U3811 ( .C1(n5809), .C2(n6741), .A(n6742), .B(n6743), .ZN(n6738) );
  aon211d1 U3812 ( .C1(n6744), .C2(n6745), .B(n6746), .A(n4191), .ZN(n6742) );
  oai22d1 U3813 ( .A1(n6748), .A2(n6741), .B1(n6749), .B2(n6750), .ZN(n6745)
         );
  aoi321d1 U3814 ( .C1(n5828), .C2(n4152), .C3(n6751), .B1(n4214), .B2(n6665), 
        .A(n4213), .ZN(n6749) );
  aoi311d1 U3815 ( .C1(n6754), .C2(n6755), .C3(n6756), .A(n6757), .B(n6758), 
        .ZN(n6751) );
  aoi21d1 U3816 ( .B1(n5042), .B2(n4153), .A(n4213), .ZN(n6758) );
  oai21d1 U3817 ( .B1(n6760), .B2(n6761), .A(n6762), .ZN(n6756) );
  aoi31d1 U3819 ( .B1(n5852), .B2(images_bus[82]), .B3(n6760), .A(n6766), .ZN(
        n6763) );
  aon211d1 U3821 ( .C1(n6770), .C2(n6771), .B(n6772), .A(n4169), .ZN(n6769) );
  oan211d1 U3822 ( .C1(images_bus[97]), .C2(n5031), .B(n6773), .A(n6774), .ZN(
        n6770) );
  aon211d1 U3823 ( .C1(n6775), .C2(n4116), .B(n4132), .A(n4064), .ZN(n6773) );
  aoi31d1 U3825 ( .B1(n6779), .B2(n5890), .B3(n6780), .A(n6781), .ZN(n6775) );
  aoi21d1 U3826 ( .B1(n5886), .B2(n6782), .A(n6783), .ZN(n6780) );
  aon211d1 U3827 ( .C1(n6784), .C2(n6785), .B(n6786), .A(n6784), .ZN(n6782) );
  aon211d1 U3828 ( .C1(n6787), .C2(n6788), .B(n6789), .A(n5895), .ZN(n6785) );
  oai321d1 U3829 ( .C1(n5905), .C2(n6790), .C3(n6791), .B1(n6792), .B2(n6791), 
        .A(n6793), .ZN(n6788) );
  aoi31d1 U3830 ( .B1(n6790), .B2(n6794), .B3(n4109), .A(n6796), .ZN(n6792) );
  aor31d1 U3833 ( .B1(n6800), .B2(n6801), .B3(n6802), .A(n6803), .Z(n6798) );
  aor311d1 U3834 ( .C1(n6802), .C2(n5921), .C3(n6804), .A(n5917), .B(n4105), 
        .Z(n6801) );
  oai211d1 U3836 ( .C1(n6809), .C2(n5017), .A(n6808), .B(n6810), .ZN(n6807) );
  oan211d1 U3837 ( .C1(n6811), .C2(n6812), .B(n4086), .A(n6814), .ZN(n6809) );
  aoi311d1 U3838 ( .C1(n6815), .C2(n6816), .C3(n4134), .A(n7603), .B(n6812), 
        .ZN(n6811) );
  oai31d1 U3840 ( .B1(n6819), .B2(n4090), .B3(n6820), .A(n6821), .ZN(n6816) );
  oan211d1 U3841 ( .C1(n6822), .C2(n6823), .B(n6824), .A(n5030), .ZN(n6820) );
  aoi211d1 U3842 ( .C1(n5024), .C2(n6825), .A(n4133), .B(n6827), .ZN(n6822) );
  oan211d1 U3843 ( .C1(n6828), .C2(n6829), .B(images_bus[121]), .A(n6830), 
        .ZN(n6827) );
  oai321d1 U3845 ( .C1(n6833), .C2(n6834), .C3(n6835), .B1(n6836), .B2(n6835), 
        .A(n5449), .ZN(n6832) );
  aon211d1 U3846 ( .C1(n3999), .C2(n6649), .B(n6839), .A(n4057), .ZN(n6833) );
  oan211d1 U3847 ( .C1(n6841), .C2(n4002), .B(n6843), .A(n5041), .ZN(n6839) );
  aoi22d1 U3848 ( .A1(n4391), .A2(n6844), .B1(n6845), .B2(n4006), .ZN(n6841)
         );
  oai21d1 U3849 ( .B1(n5055), .B2(n6846), .A(n6847), .ZN(n6844) );
  nd13d1 U3850 ( .A1(n6848), .A2(n6845), .A3(images_bus[131]), .ZN(n6847) );
  aon211d1 U3851 ( .C1(n6845), .C2(n4735), .B(n6850), .A(n6851), .ZN(n6846) );
  aoi31d1 U3853 ( .B1(n6854), .B2(n4053), .B3(n6856), .A(n6857), .ZN(n6852) );
  oai31d1 U3856 ( .B1(n6863), .B2(n7023), .B3(n5440), .A(n6864), .ZN(n6862) );
  aon211d1 U3857 ( .C1(n6865), .C2(n4043), .B(n6867), .A(n6868), .ZN(n6864) );
  aoi31d1 U3858 ( .B1(n6869), .B2(n6870), .B3(images_bus[160]), .A(n5117), 
        .ZN(n6867) );
  aon211d1 U3859 ( .C1(n3913), .C2(n6872), .B(n5762), .A(n5120), .ZN(n6869) );
  oai21d1 U3860 ( .B1(n6873), .B2(n6874), .A(n3900), .ZN(n6872) );
  aoi211d1 U3862 ( .C1(n3914), .C2(n5278), .A(n6877), .B(n6876), .ZN(n6873) );
  oai222d1 U3863 ( .A1(images_bus[165]), .A2(n6878), .B1(n6879), .B2(n6880), 
        .C1(n6881), .C2(n3915), .ZN(n6877) );
  aoi211d1 U3865 ( .C1(n3922), .C2(n5994), .A(n6885), .B(n6886), .ZN(n6879) );
  aoi31d1 U3866 ( .B1(n6881), .B2(n6887), .B3(n6888), .A(n6889), .ZN(n6886) );
  aon211d1 U3867 ( .C1(n3924), .C2(n6891), .B(n5139), .A(n3923), .ZN(n6887) );
  aon211d1 U3869 ( .C1(n3901), .C2(n6895), .B(n6896), .A(n5141), .ZN(n6891) );
  aoi31d1 U3870 ( .B1(n3929), .B2(n5189), .B3(n3927), .A(n5676), .ZN(n5141) );
  aor31d1 U3871 ( .B1(n5192), .B2(n6898), .B3(n3901), .A(n6899), .Z(n6895) );
  aon211d1 U3872 ( .C1(n3932), .C2(n6900), .B(n3931), .A(n6902), .ZN(n6898) );
  oai211d1 U3873 ( .C1(n6903), .C2(n5158), .A(n6904), .B(n6905), .ZN(n6900) );
  aon211d1 U3874 ( .C1(n6906), .C2(n6907), .B(n5949), .A(n3935), .ZN(n6904) );
  oan211d1 U3876 ( .C1(n6909), .C2(n6907), .B(n6910), .A(n5558), .ZN(n6903) );
  aoi31d1 U3877 ( .B1(n6911), .B2(n6912), .B3(n3941), .A(n6913), .ZN(n6909) );
  aon211d1 U3880 ( .C1(images_bus[183]), .C2(n6916), .B(n6917), .A(n6918), 
        .ZN(n6915) );
  aon211d1 U3881 ( .C1(n3962), .C2(n6920), .B(n6921), .A(n3952), .ZN(n6916) );
  oai211d1 U3882 ( .C1(n4958), .C2(n3959), .A(images_bus[185]), .B(n6924), 
        .ZN(n6920) );
  aoi31d1 U3884 ( .B1(n6929), .B2(n4958), .B3(n6928), .A(n6930), .ZN(n6925) );
  aon211d1 U3885 ( .C1(n3956), .C2(n6932), .B(n5769), .A(N10551), .ZN(n6929)
         );
  oai221d1 U3886 ( .B1(n6933), .B2(n3818), .C1(n6627), .C2(n5193), .A(
        images_bus[189]), .ZN(n6932) );
  aoi31d1 U3889 ( .B1(n6937), .B2(n3882), .B3(n6939), .A(n6940), .ZN(n6933) );
  oan211d1 U3891 ( .C1(n6943), .C2(n6944), .B(n6945), .A(n6016), .ZN(n6937) );
  aon211d1 U3892 ( .C1(n3890), .C2(images_bus[204]), .B(n6947), .A(n3840), 
        .ZN(n6945) );
  oan211d1 U3895 ( .C1(n5548), .C2(n3891), .B(n6954), .A(n3846), .ZN(n6952) );
  aon211d1 U3897 ( .C1(n6956), .C2(n6957), .B(n6958), .A(n3851), .ZN(n6954) );
  oan211d1 U3899 ( .C1(n6962), .C2(n6963), .B(n3862), .A(n6964), .ZN(n6959) );
  oan211d1 U3901 ( .C1(n6968), .C2(n5747), .B(n6969), .A(n6970), .ZN(n6965) );
  aoi31d1 U3902 ( .B1(n6971), .B2(n6972), .B3(n6973), .A(n5279), .ZN(n6968) );
  oai211d1 U3903 ( .C1(n6974), .C2(n3746), .A(n6976), .B(n3740), .ZN(n6972) );
  aoi31d1 U3905 ( .B1(n3748), .B2(n6025), .B3(n3757), .A(n4691), .ZN(n5290) );
  oan211d1 U3906 ( .C1(n6977), .C2(n6978), .B(n3621), .A(n5289), .ZN(n6974) );
  aoi311d1 U3908 ( .C1(n6981), .C2(n7153), .C3(n3807), .A(n6980), .B(n5296), 
        .ZN(n6977) );
  oai222d1 U3909 ( .A1(n6983), .A2(n4407), .B1(n6984), .B2(n4407), .C1(
        images_bus[233]), .C2(n6985), .ZN(n6981) );
  aoim31d1 U3910 ( .B1(n6986), .B2(n6987), .B3(n6988), .A(n6989), .ZN(n6984)
         );
  aoi311d1 U3911 ( .C1(n3770), .C2(n6991), .C3(n3801), .A(n6992), .B(n3650), 
        .ZN(n6986) );
  oai211d1 U3913 ( .C1(n5544), .C2(n5317), .A(n6994), .B(n6995), .ZN(n6991) );
  aoi21d1 U3914 ( .B1(n3774), .B2(n6996), .A(n3771), .ZN(n6995) );
  aoi31d1 U3916 ( .B1(n3800), .B2(n5542), .B3(n3774), .A(n5937), .ZN(n5310) );
  aon211d1 U3918 ( .C1(n3777), .C2(n2803), .B(n5063), .A(n6999), .ZN(n6994) );
  aoim211d1 U3920 ( .C1(n7001), .C2(n7002), .A(n6996), .B(n5323), .ZN(n7000)
         );
  aoi211d1 U3922 ( .C1(n7005), .C2(n5331), .A(n3653), .B(n5332), .ZN(n7001) );
  aoi31d1 U3923 ( .B1(n7007), .B2(n7008), .B3(n7009), .A(n5326), .ZN(n7005) );
  oai31d1 U3925 ( .B1(n7013), .B2(n7014), .B3(n7015), .A(n3791), .ZN(n7010) );
  aoi31d1 U3926 ( .B1(n3789), .B2(n7018), .B3(n3575), .A(n7020), .ZN(n7014) );
  aoi322d1 U3928 ( .C1(n3524), .C2(n3531), .C3(n7024), .A1(n5348), .A2(n7025), 
        .B1(n7026), .B2(n7027), .ZN(n7021) );
  oan211d1 U3929 ( .C1(n7028), .C2(n7029), .B(n7030), .A(n7031), .ZN(n7024) );
  oai211d1 U3930 ( .C1(n7032), .C2(n7033), .A(n5745), .B(n3539), .ZN(n7030) );
  oai211d1 U3933 ( .C1(n7038), .C2(n7039), .A(n7040), .B(n3542), .ZN(n7036) );
  oan211d1 U3935 ( .C1(n12169), .C2(n3513), .B(n7043), .A(n7044), .ZN(n7038)
         );
  oai211d1 U3937 ( .C1(images_bus[289]), .C2(n5382), .A(n7049), .B(n3486), 
        .ZN(n7048) );
  oai31d1 U3939 ( .B1(n7052), .B2(n5738), .B3(n7051), .A(n7053), .ZN(n7049) );
  aon211d1 U3940 ( .C1(n7054), .C2(n7055), .B(n5383), .A(n7056), .ZN(n7052) );
  aon211d1 U3941 ( .C1(n3473), .C2(n5265), .B(n4483), .A(n3474), .ZN(n7056) );
  oan211d1 U3943 ( .C1(n7059), .C2(n7060), .B(n7061), .A(n3427), .ZN(n7058) );
  aon211d1 U3945 ( .C1(n3470), .C2(n7063), .B(n6007), .A(n7064), .ZN(n7060) );
  aon211d1 U3946 ( .C1(n7065), .C2(images_bus[297]), .B(n5396), .A(n6018), 
        .ZN(n7063) );
  aoi22d1 U3947 ( .A1(n3464), .A2(n7068), .B1(n3466), .B2(n7070), .ZN(n7065)
         );
  aon211d1 U3948 ( .C1(n7071), .C2(n3489), .B(n5395), .A(images_bus[299]), 
        .ZN(n7068) );
  oan211d1 U3949 ( .C1(n7073), .C2(n7074), .B(n3431), .A(n5164), .ZN(n7071) );
  aoi31d1 U3950 ( .B1(n3489), .B2(n4438), .B3(n7077), .A(n7078), .ZN(n7073) );
  aoi322d1 U3951 ( .C1(n3438), .C2(n7080), .C3(n3434), .A1(n3460), .A2(n5931), 
        .B1(n7082), .B2(n7083), .ZN(n7077) );
  oan211d1 U3952 ( .C1(n7084), .C2(n7085), .B(images_bus[305]), .A(n6183), 
        .ZN(n7083) );
  aoi321d1 U3954 ( .C1(n7088), .C2(images_bus[307]), .C3(n7089), .B1(
        images_bus[307]), .B2(n7090), .A(n5412), .ZN(n7086) );
  aoi21d1 U3955 ( .B1(n7091), .B2(n7092), .A(n3455), .ZN(n7089) );
  oai211d1 U3958 ( .C1(n3448), .C2(n7098), .A(n7099), .B(n7100), .ZN(n7096) );
  oai31d1 U3960 ( .B1(n3487), .B2(n3446), .B3(n4993), .A(n7106), .ZN(n7101) );
  aon211d1 U3963 ( .C1(n7111), .C2(n3365), .B(n7112), .A(n5424), .ZN(n7107) );
  aoi21d1 U3965 ( .B1(n7113), .B2(n7114), .A(n6197), .ZN(n7111) );
  aon211d1 U3966 ( .C1(n3355), .C2(images_bus[323]), .B(n7116), .A(n3417), 
        .ZN(n7113) );
  oan211d1 U3968 ( .C1(n7118), .C2(n4547), .B(n7119), .A(n4538), .ZN(n7116) );
  aoi311d1 U3969 ( .C1(n3410), .C2(n7120), .C3(n3409), .A(n3354), .B(n7122), 
        .ZN(n7118) );
  oai31d1 U3970 ( .B1(n7123), .B2(n7124), .B3(n7125), .A(n7126), .ZN(n7120) );
  aoi31d1 U3971 ( .B1(n3375), .B2(n7128), .B3(n7129), .A(n3354), .ZN(n7124) );
  aoi21d1 U3972 ( .B1(n7130), .B2(n7131), .A(n7132), .ZN(n7129) );
  oai211d1 U3973 ( .C1(n3353), .C2(n7134), .A(n7135), .B(n3380), .ZN(n7130) );
  oan211d1 U3975 ( .C1(n7138), .C2(n7139), .B(n7140), .A(n7141), .ZN(n7134) );
  aoi311d1 U3976 ( .C1(n7142), .C2(n3273), .C3(n7143), .A(n7144), .B(n7145), 
        .ZN(n7138) );
  aoi311d1 U3978 ( .C1(n6283), .C2(n5475), .C3(images_bus[352]), .A(n7147), 
        .B(n7148), .ZN(n7143) );
  aoi322d1 U3980 ( .C1(n2804), .C2(n7154), .C3(n3325), .A1(n7156), .A2(n7157), 
        .B1(n5720), .B2(n4586), .ZN(n7151) );
  oan211d1 U3981 ( .C1(n7158), .C2(n7159), .B(n7160), .A(n4586), .ZN(n7156) );
  oai21d1 U3984 ( .B1(n7162), .B2(n7163), .A(n7164), .ZN(n7159) );
  oai211d1 U3986 ( .C1(n7168), .C2(n7169), .A(n5626), .B(n7170), .ZN(n7167) );
  aoi31d1 U3988 ( .B1(n3257), .B2(n7174), .B3(n3280), .A(n3314), .ZN(n7172) );
  aon211d1 U3990 ( .C1(n3289), .C2(n7177), .B(n7178), .A(n6316), .ZN(n7174) );
  oai211d1 U3991 ( .C1(n7179), .C2(n7180), .A(n7181), .B(n3255), .ZN(n7177) );
  aon211d1 U3993 ( .C1(n3288), .C2(n6597), .B(n5920), .A(n3286), .ZN(n7181) );
  aoi31d1 U3995 ( .B1(n7186), .B2(n6327), .B3(n7187), .A(n5491), .ZN(n7185) );
  aoi21d1 U3998 ( .B1(n3308), .B2(n7193), .A(n3311), .ZN(n7192) );
  oai211d1 U4003 ( .C1(n5380), .C2(n7197), .A(n7198), .B(n7199), .ZN(n7196) );
  aoi21d1 U4004 ( .B1(n6342), .B2(n7200), .A(n7201), .ZN(n7199) );
  oai211d1 U4005 ( .C1(n7202), .C2(n6353), .A(images_bus[379]), .B(n7203), 
        .ZN(n7200) );
  aoi321d1 U4007 ( .C1(n3297), .C2(n3168), .C3(n7204), .B1(n3297), .B2(n3138), 
        .A(n3256), .ZN(n7202) );
  aoi31d1 U4009 ( .B1(n7206), .B2(n3161), .B3(n7208), .A(n7209), .ZN(n7204) );
  aoi211d1 U4010 ( .C1(n3167), .C2(n7210), .A(n7211), .B(n7212), .ZN(n7208) );
  aoi31d1 U4012 ( .B1(n7216), .B2(n7217), .B3(n7218), .A(n7210), .ZN(n7213) );
  aoi21d1 U4013 ( .B1(n7219), .B2(n7220), .A(n6364), .ZN(n7218) );
  aor311d1 U4014 ( .C1(n7221), .C2(n7220), .C3(n3143), .A(n7223), .B(n4655), 
        .Z(n7219) );
  aor211d1 U4015 ( .C1(n7224), .C2(n3143), .A(n7225), .B(n6380), .Z(n7221) );
  aon211d1 U4017 ( .C1(n7227), .C2(n7228), .B(n7229), .A(n7230), .ZN(n7224) );
  oai211d1 U4018 ( .C1(n7231), .C2(n3196), .A(n7233), .B(n7234), .ZN(n7228) );
  aon211d1 U4019 ( .C1(images_bus[399]), .C2(n7235), .B(n7236), .A(n7229), 
        .ZN(n7234) );
  aon211d1 U4020 ( .C1(n3207), .C2(n7238), .B(n7239), .A(n3198), .ZN(n7233) );
  oan211d1 U4022 ( .C1(n3235), .C2(n4302), .B(n3239), .A(n3144), .ZN(n7239) );
  oai322d1 U4023 ( .C1(n3144), .C2(n3211), .C3(n4302), .A1(n7246), .A2(n7247), 
        .B1(n7248), .B2(n7249), .ZN(n7238) );
  aoi31d1 U4024 ( .B1(images_bus[407]), .B2(n3211), .B3(n7250), .A(n6406), 
        .ZN(n7248) );
  aoi311d1 U4025 ( .C1(n3220), .C2(n6587), .C3(n7252), .A(n7253), .B(n7254), 
        .ZN(n7246) );
  oan211d1 U4026 ( .C1(n3228), .C2(n7256), .B(n7257), .A(n7258), .ZN(n7254) );
  oai211d1 U4028 ( .C1(n7263), .C2(n4707), .A(n4708), .B(n7264), .ZN(n7262) );
  aoi22d1 U4029 ( .A1(n4710), .A2(n3025), .B1(n7266), .B2(n4713), .ZN(n7264)
         );
  aoi211d1 U4030 ( .C1(n4715), .C2(n7267), .A(n7268), .B(n7269), .ZN(n7263) );
  aoi21d1 U4031 ( .B1(n4721), .B2(n4720), .A(n7270), .ZN(n7269) );
  oai211d1 U4032 ( .C1(n3127), .C2(n7270), .A(n7272), .B(n7273), .ZN(n7267) );
  oai21d1 U4035 ( .B1(n4731), .B2(n5583), .A(n4724), .ZN(n7277) );
  oai211d1 U4036 ( .C1(n3065), .C2(n7276), .A(n3063), .B(n7279), .ZN(n7275) );
  aoi22d1 U4037 ( .A1(n3064), .A2(n7280), .B1(n4741), .B2(n7281), .ZN(n7279)
         );
  oai21d1 U4038 ( .B1(n5703), .B2(n4739), .A(n5589), .ZN(n4741) );
  oaim22d1 U4039 ( .A1(n7282), .A2(n5597), .B1(n4744), .B2(n7281), .ZN(n7280)
         );
  aoi211d1 U4040 ( .C1(n5600), .C2(n7281), .A(n7283), .B(n7284), .ZN(n7282) );
  oai22d1 U4041 ( .A1(n5602), .A2(n7285), .B1(n7286), .B2(n3082), .ZN(n7283)
         );
  aoim2m11d1 U4043 ( .C1(n7285), .C2(n3090), .B(n7289), .A(n7290), .ZN(n7286)
         );
  oai22d1 U4044 ( .A1(n7291), .A2(n3087), .B1(n7292), .B2(n5616), .ZN(n7290)
         );
  aoi311d1 U4045 ( .C1(n2946), .C2(n7294), .C3(n7295), .A(n7296), .B(n2921), 
        .ZN(n7292) );
  aon211d1 U4047 ( .C1(n7299), .C2(n7300), .B(n7301), .A(n7302), .ZN(n7298) );
  aor21d1 U4048 ( .B1(n7303), .B2(n7304), .A(n7305), .Z(n7296) );
  oan211d1 U4049 ( .C1(n7306), .C2(n2947), .B(n7308), .A(n7309), .ZN(n7295) );
  aor311d1 U4050 ( .C1(n7310), .C2(n7311), .C3(n3004), .A(n7313), .B(n7314), 
        .Z(n7308) );
  aoi22d1 U4051 ( .A1(n7315), .A2(images_bus[457]), .B1(n7316), .B2(n7317), 
        .ZN(n7310) );
  aoi31d1 U4052 ( .B1(n3003), .B2(n7319), .B3(n7320), .A(n7321), .ZN(n7306) );
  oan211d1 U4053 ( .C1(n2928), .C2(n7323), .B(n7324), .A(n3002), .ZN(n7321) );
  aor221d1 U4056 ( .B1(n2805), .B2(n7334), .C1(n7335), .C2(images_bus[480]), 
        .A(n7336), .Z(n7330) );
  oan211d1 U4057 ( .C1(n7337), .C2(n7335), .B(n7188), .A(n7338), .ZN(n7334) );
  oai322d1 U4060 ( .C1(n7340), .C2(n7341), .C3(n2861), .A1(n7343), .A2(n7344), 
        .B1(n7345), .B2(n7346), .ZN(n7339) );
  aoi21d1 U4061 ( .B1(n2856), .B2(n7347), .A(n2854), .ZN(n7343) );
  oai211d1 U4064 ( .C1(n5696), .C2(n4876), .A(n7351), .B(n2867), .ZN(n7347) );
  aon211d1 U4066 ( .C1(n4920), .C2(n5894), .B(n7354), .A(n2874), .ZN(n7353) );
  aon211d1 U4070 ( .C1(images_bus[461]), .C2(n7359), .B(n7336), .A(
        images_bus[460]), .ZN(n7323) );
  aoi21d1 U4081 ( .B1(n3117), .B2(n7362), .A(n4749), .ZN(n5602) );
  oai221d1 U4084 ( .B1(n3065), .B2(n4950), .C1(n3070), .C2(n4739), .A(n7364), 
        .ZN(n4737) );
  oai31d1 U4092 ( .B1(n7368), .B2(n5806), .B3(n7249), .A(n7369), .ZN(n7253) );
  oai211d1 U4093 ( .C1(n6441), .C2(n7370), .A(n6430), .B(n3145), .ZN(n7369) );
  aoi211d1 U4096 ( .C1(n6084), .C2(n3128), .A(n3037), .B(n6160), .ZN(n6441) );
  aor21d1 U4099 ( .B1(n7258), .B2(n4901), .A(n7374), .Z(n6587) );
  oan211d1 U4103 ( .C1(n6736), .C2(n6401), .B(n3205), .A(n3197), .ZN(n7376) );
  oan211d1 U4116 ( .C1(n7383), .C2(n5988), .B(n3318), .A(n4653), .ZN(n7162) );
  oan211d1 U4117 ( .C1(n7384), .C2(n7385), .B(n7170), .A(n7386), .ZN(n7383) );
  aoi31d1 U4136 ( .B1(n7103), .B2(n3444), .B3(n7392), .A(n7394), .ZN(n7098) );
  aon211d1 U4141 ( .C1(n3452), .C2(n5826), .B(n7396), .A(n3454), .ZN(n7095) );
  aoi21d1 U4157 ( .B1(n3517), .B2(n7012), .A(n7409), .ZN(n7026) );
  aor31d1 U4166 ( .B1(n6962), .B2(images_bus[222]), .B3(images_bus[223]), .A(
        n7242), .Z(n6970) );
  aon211d1 U4167 ( .C1(n3809), .C2(n5754), .B(n5268), .A(n3742), .ZN(n6971) );
  aon211d1 U4179 ( .C1(n3943), .C2(n7426), .B(n7427), .A(n3939), .ZN(n6911) );
  oai21d1 U4180 ( .B1(n6918), .B2(n7428), .A(images_bus[181]), .ZN(n7426) );
  aoi21d1 U4211 ( .B1(n5957), .B2(n4108), .A(n7442), .ZN(n5921) );
  aoi21d1 U4216 ( .B1(n7444), .B2(n6772), .A(n7251), .ZN(n6779) );
  aoi311d1 U4238 ( .C1(n7459), .C2(images_bus[16]), .C3(n7460), .A(n7461), .B(
        n6678), .ZN(N26362) );
  nd13d1 U4239 ( .A1(n7462), .A2(n7463), .A3(n7464), .ZN(n6678) );
  aoi211d1 U4241 ( .C1(n7468), .C2(n7469), .A(n4580), .B(n7471), .ZN(n7460) );
  aoi22d1 U4242 ( .A1(n7472), .A2(n7473), .B1(n6681), .B2(n7474), .ZN(n7459)
         );
  oai211d1 U4243 ( .C1(n7475), .C2(n4361), .A(n7477), .B(n7478), .ZN(n7474) );
  aon211d1 U4245 ( .C1(n7483), .C2(n7484), .B(n7485), .A(n7486), .ZN(n7480) );
  aoi31d1 U4246 ( .B1(n7487), .B2(n7488), .B3(n7489), .A(n7490), .ZN(n7479) );
  oan211d1 U4247 ( .C1(n7491), .C2(n7492), .B(n7493), .A(n7494), .ZN(n7489) );
  oaim22d1 U4248 ( .A1(n7495), .A2(n7496), .B1(n4291), .B2(n7498), .ZN(n7492)
         );
  aoi31d1 U4249 ( .B1(n6691), .B2(n7499), .B3(n7500), .A(n4291), .ZN(n7495) );
  oai221d1 U4250 ( .B1(n7501), .B2(n5800), .C1(n7502), .C2(n4287), .A(n7504), 
        .ZN(n7499) );
  aoi31d1 U4252 ( .B1(images_bus[45]), .B2(images_bus[44]), .B3(n7505), .A(
        n7506), .ZN(n7501) );
  aoi31d1 U4253 ( .B1(n7507), .B2(n7508), .B3(n7509), .A(n4251), .ZN(n7506) );
  aoi211d1 U4254 ( .C1(n7511), .C2(n7512), .A(n7513), .B(n4288), .ZN(n7509) );
  aoi21d1 U4256 ( .B1(n6727), .B2(n7516), .A(n4257), .ZN(n7508) );
  oai211d1 U4258 ( .C1(n7518), .C2(n6730), .A(n4263), .B(n4290), .ZN(n7516) );
  aoi31d1 U4261 ( .B1(n4289), .B2(n4205), .B3(n7526), .A(n7527), .ZN(n7523) );
  aoi22d1 U4262 ( .A1(n7528), .A2(n7529), .B1(n7530), .B2(n4210), .ZN(n7526)
         );
  oan211d1 U4263 ( .C1(n6403), .C2(n7532), .B(n7533), .A(n7534), .ZN(n7528) );
  oai311d1 U4264 ( .C1(n7535), .C2(n7536), .C3(n7537), .A(n4152), .B(n4149), 
        .ZN(n7533) );
  aon211d1 U4266 ( .C1(n4209), .C2(images_bus[76]), .B(n7543), .A(
        images_bus[77]), .ZN(n7540) );
  aoi31d1 U4267 ( .B1(n7544), .B2(n7545), .B3(n7546), .A(n6667), .ZN(n7543) );
  oai21d1 U4268 ( .B1(n5842), .B2(n7547), .A(n7548), .ZN(n7546) );
  aon211d1 U4269 ( .C1(n4173), .C2(n7550), .B(n7551), .A(n5023), .ZN(n7544) );
  aoi221d1 U4271 ( .B1(n7556), .B2(n7557), .C1(n4160), .C2(n7559), .A(n5106), 
        .ZN(n7555) );
  oan211d1 U4272 ( .C1(n7560), .C2(n7561), .B(n7562), .A(n5861), .ZN(n7556) );
  aoi22d1 U4273 ( .A1(n4166), .A2(n7563), .B1(N9106), .B2(n5456), .ZN(n7560)
         );
  oan211d1 U4276 ( .C1(n7569), .C2(n7570), .B(n7571), .A(n7572), .ZN(n7568) );
  nd13d1 U4277 ( .A1(n7573), .A2(n4110), .A3(n7575), .ZN(n7571) );
  oan211d1 U4278 ( .C1(n5917), .C2(n7576), .B(n7577), .A(n7578), .ZN(n7575) );
  aon211d1 U4279 ( .C1(n4108), .C2(n7579), .B(n7580), .A(n5914), .ZN(n7576) );
  oai322d1 U4280 ( .C1(n7581), .C2(n7582), .C3(n7583), .A1(n7584), .A2(n7585), 
        .B1(n4083), .B2(n7581), .ZN(n7579) );
  ora211d1 U4281 ( .C1(n5017), .C2(n7587), .A(n7584), .B(n6810), .Z(n7582) );
  aoi21d1 U4282 ( .B1(n4082), .B2(n4084), .A(n5575), .ZN(n6810) );
  ora211d1 U4284 ( .C1(n7589), .C2(n7590), .A(n5579), .B(n7584), .Z(n7587) );
  oan211d1 U4285 ( .C1(n7591), .C2(n7592), .B(n6821), .A(n4101), .ZN(n7589) );
  oan211d1 U4287 ( .C1(n5030), .C2(n7593), .B(n7439), .A(n7594), .ZN(n7591) );
  oai22d1 U4288 ( .A1(n7595), .A2(n7596), .B1(n7596), .B2(n7597), .ZN(n7593)
         );
  aon211d1 U4289 ( .C1(n5449), .C2(n7598), .B(n7599), .A(n7600), .ZN(n7597) );
  aoi31d1 U4291 ( .B1(n7600), .B2(n6831), .B3(n7601), .A(n6830), .ZN(n7595) );
  oan211d1 U4292 ( .C1(n7602), .C2(n4129), .B(n4097), .A(n6825), .ZN(n7601) );
  aoi311d1 U4294 ( .C1(n3995), .C2(n7607), .C3(n7605), .A(n6834), .B(n5951), 
        .ZN(n7602) );
  aon211d1 U4295 ( .C1(n7608), .C2(n7609), .B(n7610), .A(n4000), .ZN(n7607) );
  oan211d1 U4296 ( .C1(n3989), .C2(n5054), .B(n7613), .A(n5768), .ZN(n7608) );
  aoi211d1 U4298 ( .C1(n7617), .C2(n7618), .A(n5050), .B(n7619), .ZN(n7616) );
  oai211d1 U4300 ( .C1(n7623), .C2(n5084), .A(n7624), .B(n4030), .ZN(n7622) );
  aoi211d1 U4302 ( .C1(n5088), .C2(n7627), .A(n7628), .B(n5090), .ZN(n7623) );
  aon211d1 U4303 ( .C1(n7629), .C2(n7630), .B(n7631), .A(n5101), .ZN(n7627) );
  aoi221d1 U4304 ( .B1(n4035), .B2(n7023), .C1(n7633), .C2(n7634), .A(n7635), 
        .ZN(n7630) );
  aon211d1 U4306 ( .C1(n4042), .C2(n7640), .B(n5103), .A(n4033), .ZN(n7638) );
  oai31d1 U4307 ( .B1(n7642), .B2(n7643), .B3(n3907), .A(n4032), .ZN(n7637) );
  ora311d1 U4309 ( .C1(n7645), .C2(n7646), .C3(n7642), .A(n7647), .B(n7648), 
        .Z(n7643) );
  aoim21d1 U4310 ( .B1(n7649), .B2(n6123), .A(n7650), .ZN(n7646) );
  aoi31d1 U4312 ( .B1(n7654), .B2(n5163), .B3(n7655), .A(n3976), .ZN(n7651) );
  aoi31d1 U4314 ( .B1(n7658), .B2(n7659), .B3(n7660), .A(n5144), .ZN(n7655) );
  oai31d1 U4315 ( .B1(n7661), .B2(n7662), .B3(n6914), .A(n3937), .ZN(n7658) );
  aoi31d1 U4316 ( .B1(n3977), .B2(n7665), .B3(n7666), .A(n7667), .ZN(n7662) );
  oai311d1 U4317 ( .C1(n7668), .C2(n7661), .C3(n7669), .A(n3953), .B(n6003), 
        .ZN(n7665) );
  oai21d1 U4318 ( .B1(n7670), .B2(n6632), .A(n7671), .ZN(n7668) );
  oai22d1 U4321 ( .A1(n7675), .A2(n7676), .B1(n4402), .B2(n7677), .ZN(n7672)
         );
  aon211d1 U4322 ( .C1(n3887), .C2(n3841), .B(n7680), .A(n3845), .ZN(n7677) );
  oai21d1 U4323 ( .B1(n7682), .B2(n5215), .A(n7683), .ZN(n7680) );
  aoi31d1 U4325 ( .B1(images_bus[205]), .B2(images_bus[204]), .B3(n3887), .A(
        n7686), .ZN(n7682) );
  aoi31d1 U4326 ( .B1(n3847), .B2(n7688), .B3(n7689), .A(n7690), .ZN(n7686) );
  aoi31d1 U4327 ( .B1(n7691), .B2(n7692), .B3(n6046), .A(n7693), .ZN(n7689) );
  aon211d1 U4329 ( .C1(n7695), .C2(n7696), .B(n7079), .A(n7697), .ZN(n7688) );
  aoi31d1 U4330 ( .B1(n3888), .B2(n6052), .B3(n7699), .A(n7700), .ZN(n7695) );
  aoi22d1 U4331 ( .A1(n3867), .A2(n7702), .B1(n3866), .B2(n7704), .ZN(n7699)
         );
  aon211d1 U4333 ( .C1(n7708), .C2(n7709), .B(n7710), .A(n6055), .ZN(n7707) );
  aon211d1 U4334 ( .C1(n3721), .C2(n7711), .B(n7712), .A(n6053), .ZN(n7706) );
  oan211d1 U4335 ( .C1(n7713), .C2(n5287), .B(n7714), .A(n4425), .ZN(n7712) );
  oan211d1 U4337 ( .C1(n7714), .C2(n7716), .B(n7717), .A(n5286), .ZN(n7715) );
  oai22d1 U4339 ( .A1(n6987), .A2(n7721), .B1(n7722), .B2(n3803), .ZN(n7720)
         );
  oan211d1 U4341 ( .C1(n7725), .C2(n7726), .B(n3769), .A(n7728), .ZN(n7722) );
  aon211d1 U4343 ( .C1(n3779), .C2(n7729), .B(n7730), .A(n3775), .ZN(n7726) );
  oan211d1 U4344 ( .C1(n7732), .C2(n7733), .B(n3776), .A(n7725), .ZN(n7730) );
  oan211d1 U4346 ( .C1(n6103), .C2(n6105), .B(n7736), .A(n6106), .ZN(n7735) );
  aor211d1 U4347 ( .C1(n7737), .C2(n3782), .A(n5750), .B(n6105), .Z(n7733) );
  oai21d1 U4348 ( .B1(n7011), .B2(n7739), .A(n7007), .ZN(n7737) );
  oai211d1 U4350 ( .C1(n7741), .C2(n7742), .A(n7743), .B(n3783), .ZN(n7732) );
  aoi221d1 U4351 ( .B1(n3572), .B2(n7746), .C1(n3521), .C2(n5350), .A(n6620), 
        .ZN(n7741) );
  oaim211d1 U4353 ( .C1(n7748), .C2(n5348), .A(n7749), .B(n5345), .ZN(n7746)
         );
  aon211d1 U4354 ( .C1(n4683), .C2(n7748), .B(n7750), .A(n3523), .ZN(n7749) );
  oan211d1 U4357 ( .C1(n7754), .C2(n7755), .B(n7756), .A(n6128), .ZN(n7750) );
  oai211d1 U4358 ( .C1(n7757), .C2(n7758), .A(n5745), .B(n7759), .ZN(n7756) );
  oan211d1 U4360 ( .C1(n7761), .C2(n7762), .B(n7763), .A(n7764), .ZN(n7757) );
  oai21d1 U4361 ( .B1(n7765), .B2(n7766), .A(n3560), .ZN(n7763) );
  aoi31d1 U4362 ( .B1(n7761), .B2(n4461), .B3(n7768), .A(n7041), .ZN(n7765) );
  aoi22d1 U4363 ( .A1(n4466), .A2(n7769), .B1(n4468), .B2(n7770), .ZN(n7768)
         );
  oai211d1 U4364 ( .C1(n3514), .C2(n3551), .A(n7772), .B(n4473), .ZN(n7770) );
  oai31d1 U4365 ( .B1(n7773), .B2(n7774), .B3(n7769), .A(n4476), .ZN(n7772) );
  oaim22d1 U4366 ( .A1(n7775), .A2(n7776), .B1(n7777), .B2(n3425), .ZN(n7773)
         );
  aoi31d1 U4367 ( .B1(n3467), .B2(n7780), .B3(n3429), .A(n7782), .ZN(n7775) );
  oai22d1 U4369 ( .A1(n7078), .A2(n7784), .B1(n7785), .B2(n7786), .ZN(n7780)
         );
  aoi221d1 U4370 ( .B1(n3437), .B2(n5531), .C1(n3438), .C2(n7072), .A(n7788), 
        .ZN(n7785) );
  aoi31d1 U4371 ( .B1(n7789), .B2(n7790), .B3(n7791), .A(n5403), .ZN(n7788) );
  aon211d1 U4372 ( .C1(n7792), .C2(n7396), .B(n7793), .A(n3457), .ZN(n7790) );
  aoi31d1 U4373 ( .B1(n7791), .B2(n5731), .B3(n7795), .A(n7796), .ZN(n7793) );
  aoi211d1 U4374 ( .C1(n7797), .C2(n7798), .A(n7799), .B(n7800), .ZN(n7795) );
  aoi31d1 U4375 ( .B1(n3499), .B2(images_bus[313]), .B3(n7802), .A(n7803), 
        .ZN(n7800) );
  aoi221d1 U4376 ( .B1(n7804), .B2(n6604), .C1(n3440), .C2(n7806), .A(n7807), 
        .ZN(n7802) );
  oai311d1 U4377 ( .C1(n6198), .C2(images_bus[319]), .C3(n6188), .A(n7808), 
        .B(n7809), .ZN(n7806) );
  aoi311d1 U4378 ( .C1(n4522), .C2(n4528), .C3(n7810), .A(n7811), .B(n7812), 
        .ZN(n7809) );
  aoim21d1 U4379 ( .B1(n7813), .B2(n7814), .A(n4536), .ZN(n7810) );
  oan211d1 U4380 ( .C1(n7815), .C2(n6215), .B(n7816), .A(n7817), .ZN(n7813) );
  aon211d1 U4381 ( .C1(n7818), .C2(n2797), .B(n7820), .A(n3414), .ZN(n7815) );
  aon211d1 U4383 ( .C1(n7823), .C2(n7824), .B(n7820), .A(n3410), .ZN(n7822) );
  aon211d1 U4384 ( .C1(n7825), .C2(n7826), .B(n6237), .A(n7827), .ZN(n7824) );
  aoi211d1 U4385 ( .C1(n3379), .C2(n7828), .A(n4563), .B(n6241), .ZN(n7826) );
  aoi211d1 U4386 ( .C1(n4559), .C2(n7829), .A(n7830), .B(n7831), .ZN(n7825) );
  oai211d1 U4387 ( .C1(n7832), .C2(n7833), .A(n3339), .B(n2798), .ZN(n7829) );
  oai21d1 U4389 ( .B1(n4565), .B2(n7837), .A(n4566), .ZN(n7836) );
  nd13d1 U4391 ( .A1(n7841), .A2(n7842), .A3(n3385), .ZN(n7840) );
  aon211d1 U4392 ( .C1(n3271), .C2(n7844), .B(n7845), .A(n7846), .ZN(n7839) );
  aon211d1 U4393 ( .C1(n7847), .C2(n7848), .B(n3274), .A(n7849), .ZN(n7844) );
  aon211d1 U4395 ( .C1(n3321), .C2(n7852), .B(n7853), .A(n6292), .ZN(n7847) );
  oaim2m11d1 U4396 ( .C1(n7165), .C2(n7854), .B(n7853), .A(n7855), .ZN(n7852)
         );
  oan211d1 U4397 ( .C1(n7169), .C2(n7856), .B(n7855), .A(n7857), .ZN(n7854) );
  oan211d1 U4398 ( .C1(n7858), .C2(n2799), .B(n5486), .A(n7860), .ZN(n7856) );
  oan211d1 U4400 ( .C1(n7862), .C2(n4620), .B(n3284), .A(n7860), .ZN(n7861) );
  aoi311d1 U4401 ( .C1(n7864), .C2(n4621), .C3(n7865), .A(n7866), .B(n4623), 
        .ZN(n7862) );
  aoi21d1 U4402 ( .B1(n7867), .B2(n4624), .A(n7868), .ZN(n7865) );
  aoi31d1 U4403 ( .B1(n3267), .B2(n4627), .B3(n7870), .A(n4630), .ZN(n7868) );
  aoi221d1 U4404 ( .B1(n4631), .B2(n7871), .C1(n3299), .C2(n7872), .A(n7873), 
        .ZN(n7870) );
  oan211d1 U4405 ( .C1(n3176), .C2(n7875), .B(n7876), .A(n4971), .ZN(n7873) );
  aon211d1 U4406 ( .C1(n7877), .C2(n7878), .B(n3153), .A(n3179), .ZN(n7875) );
  oai311d1 U4408 ( .C1(n7882), .C2(n7883), .C3(n7884), .A(n7881), .B(n3154), 
        .ZN(n7878) );
  aoi31d1 U4410 ( .B1(n3185), .B2(n7888), .B3(n7889), .A(n7886), .ZN(n7883) );
  oai321d1 U4411 ( .C1(n7890), .C2(n3156), .C3(n7236), .B1(n7892), .B2(n7893), 
        .A(n7894), .ZN(n7888) );
  aoi221d1 U4412 ( .B1(n4678), .B2(n7895), .C1(n4680), .C2(n7896), .A(n4682), 
        .ZN(n7892) );
  oai221d1 U4413 ( .B1(n3209), .B2(n7898), .C1(n5518), .C2(n5541), .A(n7899), 
        .ZN(n4682) );
  oai21d1 U4415 ( .B1(n5035), .B2(n7900), .A(n3210), .ZN(n5545) );
  aoim21d1 U4418 ( .B1(n7900), .B2(n7898), .A(n7902), .ZN(n5541) );
  oai211d1 U4419 ( .C1(n3231), .C2(n7903), .A(n4685), .B(n7904), .ZN(n7895) );
  aoi221d1 U4420 ( .B1(n7905), .B2(n4687), .C1(n3215), .C2(n7906), .A(n3230), 
        .ZN(n7904) );
  oai211d1 U4422 ( .C1(n3227), .C2(n3155), .A(n4694), .B(n7909), .ZN(n7906) );
  aoi322d1 U4423 ( .C1(n3044), .C2(n7911), .C3(n3028), .A1(n7912), .A2(n4696), 
        .B1(n3029), .B2(n7913), .ZN(n7909) );
  oai322d1 U4424 ( .C1(n6440), .C2(n3128), .C3(n7914), .A1(n7915), .A2(n7916), 
        .B1(images_bus[413]), .B2(n3035), .ZN(n7913) );
  aon211d1 U4425 ( .C1(images_bus[416]), .C2(n7918), .B(n7919), .A(n7920), 
        .ZN(n7916) );
  aon211d1 U4428 ( .C1(n7922), .C2(n7923), .B(n7924), .A(n7925), .ZN(n7911) );
  oai211d1 U4429 ( .C1(n7926), .C2(n7927), .A(n7922), .B(n3045), .ZN(n7925) );
  aoi21d1 U4430 ( .B1(n7929), .B2(n7930), .A(n3046), .ZN(n7927) );
  aoi31d1 U4431 ( .B1(images_bus[423]), .B2(n7931), .B3(n7932), .A(n7933), 
        .ZN(n7930) );
  aon211d1 U4434 ( .C1(n3125), .C2(n7938), .B(n5617), .A(n7939), .ZN(n6454) );
  oai21d1 U4436 ( .B1(n3060), .B2(n5583), .A(n3061), .ZN(n7931) );
  aoi31d1 U4437 ( .B1(n3123), .B2(n7943), .B3(n7274), .A(n7944), .ZN(n7929) );
  aoi22d1 U4439 ( .A1(n4646), .A2(n7948), .B1(images_bus[421]), .B2(n4729), 
        .ZN(n7946) );
  oai22d1 U4440 ( .A1(n7949), .A2(n7950), .B1(n7936), .B2(n7951), .ZN(n7943)
         );
  aon211d1 U4441 ( .C1(images_bus[427]), .C2(n7952), .B(n7953), .A(n5621), 
        .ZN(n7951) );
  aoi322d1 U4445 ( .C1(n7955), .C2(n5494), .C3(n7956), .A1(n7957), .A2(n12119), 
        .B1(n3117), .B2(n7958), .ZN(n7949) );
  oai211d1 U4446 ( .C1(n7959), .C2(n4756), .A(n7960), .B(n3085), .ZN(n7958) );
  oai21d1 U4448 ( .B1(n5495), .B2(n3086), .A(n7962), .ZN(n5599) );
  oai21d1 U4449 ( .B1(n7362), .B2(n7963), .A(n12119), .ZN(n7960) );
  aoi211d1 U4450 ( .C1(n5610), .C2(n5700), .A(n7964), .B(n7965), .ZN(n7959) );
  aoi31d1 U4451 ( .B1(n7966), .B2(n7967), .B3(n7968), .A(n5616), .ZN(n7965) );
  aoi21d1 U4452 ( .B1(n7304), .B2(n5699), .A(n7305), .ZN(n7968) );
  oai22d1 U4453 ( .A1(n2919), .A2(n3099), .B1(n7970), .B2(n7971), .ZN(n7305)
         );
  oaim21d1 U4456 ( .B1(n7974), .B2(n4777), .A(n7975), .ZN(n5620) );
  oai21d1 U4458 ( .B1(n2927), .B2(n7970), .A(n5614), .ZN(n7304) );
  aoi21d1 U4459 ( .B1(n5619), .B2(n4777), .A(n7976), .ZN(n5614) );
  aoi221d1 U4462 ( .B1(n4821), .B2(n7057), .C1(n2962), .C2(n7981), .A(n7982), 
        .ZN(n7979) );
  oai211d1 U4463 ( .C1(n7983), .C2(n4837), .A(n4937), .B(n7984), .ZN(n7981) );
  aoi21d1 U4464 ( .B1(n4830), .B2(n7985), .A(n7986), .ZN(n7984) );
  aoi22d1 U4465 ( .A1(n7987), .A2(n7988), .B1(n4839), .B2(n7985), .ZN(n7983)
         );
  oai211d1 U4466 ( .C1(n7989), .C2(n4848), .A(n7990), .B(n7991), .ZN(n7988) );
  oan211d1 U4467 ( .C1(n4935), .C2(n7992), .B(n4933), .A(n7993), .ZN(n7991) );
  aoi31d1 U4468 ( .B1(n7994), .B2(n7995), .B3(n7996), .A(n4846), .ZN(n7993) );
  oai21d1 U4471 ( .B1(n2842), .B2(n4929), .A(n4857), .ZN(n7997) );
  oai211d1 U4474 ( .C1(n8007), .C2(n8008), .A(n8009), .B(n8010), .ZN(n7354) );
  aoi22d1 U4475 ( .A1(n4888), .A2(n4919), .B1(n4920), .B2(n7050), .ZN(n8010)
         );
  aoim211d1 U4478 ( .C1(n4909), .C2(n8015), .A(n8016), .B(n2891), .ZN(n8012)
         );
  oan211d1 U4479 ( .C1(n2895), .C2(n8018), .B(n8019), .A(n4904), .ZN(n8015) );
  aon211d1 U4480 ( .C1(n8020), .C2(n8021), .B(n4911), .A(n2893), .ZN(n8019) );
  oai222d1 U4482 ( .A1(n5482), .A2(n8026), .B1(n4917), .B2(n4891), .C1(n4917), 
        .C2(n8027), .ZN(n8011) );
  aon211d1 U4486 ( .C1(n7300), .C2(n7299), .B(n7301), .A(n8033), .ZN(n7966) );
  oai21d1 U4488 ( .B1(n2939), .B2(n5727), .A(n8036), .ZN(n8034) );
  oai211d1 U4489 ( .C1(n8037), .C2(n8038), .A(n2939), .B(n8039), .ZN(n8036) );
  oai211d1 U4492 ( .C1(n8042), .C2(n8043), .A(n2940), .B(n8045), .ZN(n8040) );
  oan211d1 U4493 ( .C1(n2950), .C2(n5979), .B(n8047), .A(n6358), .ZN(n8042) );
  oai21d1 U4498 ( .B1(n7062), .B2(n3090), .A(n7289), .ZN(n7964) );
  aoi21d1 U4499 ( .B1(n4772), .B2(n3089), .A(n4759), .ZN(n7289) );
  oai21d1 U4500 ( .B1(n3090), .B2(n5701), .A(n8052), .ZN(n4759) );
  oai21d1 U4503 ( .B1(n4770), .B2(n4763), .A(n4761), .ZN(n5610) );
  oan211d1 U4505 ( .C1(n7366), .C2(n4720), .B(n8055), .A(n7945), .ZN(n7926) );
  oai21d1 U4515 ( .B1(n6583), .B2(n8057), .A(n8058), .ZN(n4687) );
  oai21d1 U4520 ( .B1(n5906), .B2(n7894), .A(images_bus[400]), .ZN(n7896) );
  aor211d1 U4527 ( .C1(n8060), .C2(n8062), .A(n8063), .B(n8064), .Z(n7872) );
  aoim211d1 U4532 ( .C1(n8065), .C2(n8066), .A(n8067), .B(n5043), .ZN(n4621)
         );
  oai22d1 U4533 ( .A1(n4613), .A2(n7864), .B1(n4617), .B2(n8068), .ZN(n7858)
         );
  aoi31d1 U4536 ( .B1(n7860), .B2(images_bus[364]), .B3(n8070), .A(n7067), 
        .ZN(n8068) );
  oai21d1 U4549 ( .B1(n5927), .B2(n7827), .A(images_bus[336]), .ZN(n7830) );
  aoi31d1 U4553 ( .B1(n3345), .B2(images_bus[319]), .B3(n7808), .A(n8074), 
        .ZN(n7814) );
  aoim21d1 U4558 ( .B1(n5931), .B2(n7784), .A(n5535), .ZN(n7791) );
  aoi21d1 U4565 ( .B1(images_bus[271]), .B2(n7758), .A(n7075), .ZN(n7761) );
  oai31d1 U4572 ( .B1(n8078), .B2(n6567), .B3(n7721), .A(images_bus[240]), 
        .ZN(n7725) );
  oai311d1 U4576 ( .C1(n7709), .C2(n6115), .C3(n7711), .A(images_bus[224]), 
        .B(n5748), .ZN(n7714) );
  oai211d1 U4581 ( .C1(n7419), .C2(n7694), .A(images_bus[208]), .B(n5759), 
        .ZN(n7692) );
  aoi311d1 U4590 ( .C1(n3819), .C2(n8086), .C3(n3957), .A(n3813), .B(n4318), 
        .ZN(n7670) );
  aoim31d1 U4595 ( .B1(n7657), .B2(n7433), .B3(n8091), .A(n7081), .ZN(n7660)
         );
  oai211d1 U4596 ( .C1(n3982), .C2(n7642), .A(n5780), .B(n8092), .ZN(n7657) );
  aoi211d1 U4601 ( .C1(n8095), .C2(n8096), .A(n7628), .B(n8097), .ZN(n7629) );
  nd13d1 U4603 ( .A1(n7617), .A2(n4471), .A3(images_bus[140]), .ZN(n7624) );
  or03d0 U4611 ( .A1(n7592), .A2(n7034), .A3(n5855), .Z(n7596) );
  aoi21d1 U4613 ( .B1(images_bus[111]), .B2(n7580), .A(n7097), .ZN(n7584) );
  aon211d1 U4620 ( .C1(n8105), .C2(n8106), .B(n8107), .A(n8104), .ZN(n7565) );
  oaim21d1 U4621 ( .B1(n8103), .B2(n4117), .A(n5875), .ZN(n8106) );
  oai21d1 U4628 ( .B1(n5958), .B2(n7545), .A(images_bus[80]), .ZN(n7547) );
  oai211d1 U4635 ( .C1(n7452), .C2(n8113), .A(n5778), .B(n6666), .ZN(n7532) );
  aon211d1 U4637 ( .C1(n4216), .C2(n8115), .B(n8116), .A(n8117), .ZN(n7521) );
  aoi21d1 U4638 ( .B1(n6734), .B2(n8113), .A(n4265), .ZN(n8117) );
  aoi22d1 U4642 ( .A1(n7454), .A2(n7522), .B1(n6721), .B2(n7512), .ZN(n7507)
         );
  aoi31d1 U4645 ( .B1(n7505), .B2(images_bus[44]), .B3(n6719), .A(n7105), .ZN(
        n7515) );
  oai21d1 U4650 ( .B1(n6146), .B2(n7491), .A(n6688), .ZN(n8121) );
  aon211d1 U4651 ( .C1(n4296), .C2(n7491), .B(n8123), .A(n4374), .ZN(n7488) );
  aoi211d1 U4657 ( .C1(n8131), .C2(n8132), .A(n7184), .B(n8133), .ZN(n8128) );
  aoi31d1 U4658 ( .B1(n8134), .B2(n8135), .B3(n5705), .A(n8137), .ZN(n8133) );
  aon211d1 U4659 ( .C1(n4793), .C2(n5220), .B(n8139), .A(n4789), .ZN(n8135) );
  oai21d1 U4660 ( .B1(n8141), .B2(n8142), .A(n4776), .ZN(n8134) );
  aon211d1 U4662 ( .C1(images_bus[13]), .C2(n8145), .B(n8146), .A(
        images_bus[12]), .ZN(n8142) );
  aon211d1 U4663 ( .C1(n8147), .C2(n8148), .B(n4523), .A(n4628), .ZN(n8145) );
  oai211d1 U4664 ( .C1(images_bus[15]), .C2(n8151), .A(n8152), .B(n8153), .ZN(
        n8148) );
  oai211d1 U4665 ( .C1(n8154), .C2(n4338), .A(n4595), .B(n6681), .ZN(n8152) );
  oan211d1 U4667 ( .C1(n8158), .C2(n6679), .B(n8157), .A(n8159), .ZN(n8154) );
  oan211d1 U4668 ( .C1(n8160), .C2(n5466), .B(n8161), .A(n8162), .ZN(n8158) );
  aoi31d1 U4669 ( .B1(n4339), .B2(n7487), .B3(n8164), .A(n8165), .ZN(n8160) );
  aoi31d1 U4670 ( .B1(n4383), .B2(n8167), .B3(n4384), .A(n8168), .ZN(n8164) );
  aon211d1 U4671 ( .C1(n8169), .C2(n8170), .B(n8171), .A(images_bus[27]), .ZN(
        n8167) );
  oan211d1 U4672 ( .C1(n8172), .C2(n8173), .B(n8174), .A(n4226), .ZN(n8169) );
  oai22d1 U4674 ( .A1(n8177), .A2(n8178), .B1(n8179), .B2(n8180), .ZN(n8173)
         );
  aon211d1 U4675 ( .C1(n5784), .C2(n4286), .B(n8183), .A(n4230), .ZN(n8180) );
  oan211d1 U4678 ( .C1(n8186), .C2(n8187), .B(n8188), .A(n8187), .ZN(n8185) );
  oan211d1 U4679 ( .C1(n8189), .C2(n6711), .B(images_bus[41]), .A(n8190), .ZN(
        n8186) );
  oan211d1 U4680 ( .C1(n5205), .C2(n8191), .B(n4273), .A(n6884), .ZN(n8189) );
  oai22d1 U4681 ( .A1(n8193), .A2(n8194), .B1(n8195), .B2(n8196), .ZN(n8191)
         );
  aon211d1 U4682 ( .C1(n8197), .C2(n8198), .B(n4512), .A(n4248), .ZN(n8196) );
  aon211d1 U4684 ( .C1(n4271), .C2(n8203), .B(n8204), .A(n4250), .ZN(n8201) );
  oan211d1 U4686 ( .C1(n8207), .C2(n8208), .B(n8209), .A(n4251), .ZN(n8206) );
  aoi22d1 U4688 ( .A1(n8203), .A2(n4270), .B1(n8211), .B2(n8212), .ZN(n8209)
         );
  oai211d1 U4691 ( .C1(n8219), .C2(n6730), .A(n8220), .B(n8221), .ZN(n8218) );
  aoi211d1 U4692 ( .C1(n6734), .C2(n8222), .A(n8223), .B(n8224), .ZN(n8219) );
  aon211d1 U4693 ( .C1(n8225), .C2(n8226), .B(n8116), .A(n8227), .ZN(n8223) );
  aoi221d1 U4694 ( .B1(n8228), .B2(n8229), .C1(n4224), .C2(n4217), .A(n4203), 
        .ZN(n8226) );
  oai211d1 U4697 ( .C1(n8234), .C2(n8235), .A(images_bus[63]), .B(n8233), .ZN(
        n8229) );
  aoi31d1 U4698 ( .B1(n4189), .B2(n8237), .B3(n7529), .A(n8238), .ZN(n8234) );
  oai321d1 U4700 ( .C1(n8240), .C2(n8241), .C3(n5020), .B1(n4147), .B2(n8243), 
        .A(n8244), .ZN(n8237) );
  aon211d1 U4702 ( .C1(n4152), .C2(n8245), .B(n8246), .A(images_bus[73]), .ZN(
        n8240) );
  oai31d1 U4704 ( .B1(n8250), .B2(n8251), .B3(n8252), .A(n4153), .ZN(n8248) );
  aoi31d1 U4705 ( .B1(n4219), .B2(n4510), .B3(n8254), .A(n4155), .ZN(n8252) );
  aoi21d1 U4706 ( .B1(n4178), .B2(n5958), .A(n8257), .ZN(n8254) );
  aon211d1 U4708 ( .C1(n4171), .C2(n4218), .B(n8261), .A(n4179), .ZN(n8258) );
  aoi31d1 U4709 ( .B1(n5868), .B2(n8263), .B3(n8264), .A(n4164), .ZN(n8261) );
  oai211d1 U4711 ( .C1(n8267), .C2(n8107), .A(n8268), .B(n5872), .ZN(n8263) );
  aoi21d1 U4712 ( .B1(n5875), .B2(n8269), .A(n5027), .ZN(n8267) );
  aon211d1 U4713 ( .C1(n4062), .C2(n8271), .B(n8272), .A(n4117), .ZN(n8269) );
  oai322d1 U4714 ( .C1(n5775), .C2(n4125), .C3(n7251), .A1(n8274), .A2(n5019), 
        .B1(n7569), .B2(n8275), .ZN(n8271) );
  aoi31d1 U4715 ( .B1(images_bus[101]), .B2(n5293), .B3(n4128), .A(n8277), 
        .ZN(n8274) );
  aoi21d1 U4716 ( .B1(n4126), .B2(n8279), .A(n5032), .ZN(n8277) );
  oai211d1 U4717 ( .C1(n8280), .C2(n8281), .A(n8282), .B(images_bus[104]), 
        .ZN(n8279) );
  oai21d1 U4718 ( .B1(images_bus[105]), .B2(n5905), .A(n4126), .ZN(n8281) );
  aon211d1 U4719 ( .C1(n8283), .C2(n8284), .B(n5028), .A(n8285), .ZN(n8280) );
  oai21d1 U4720 ( .B1(n4074), .B2(n7443), .A(n4110), .ZN(n8285) );
  oai21d1 U4721 ( .B1(n8287), .B2(n4493), .A(n4079), .ZN(n8284) );
  aoi31d1 U4722 ( .B1(images_bus[109]), .B2(n8289), .B3(n8283), .A(n8290), 
        .ZN(n8287) );
  oai311d1 U4723 ( .C1(n4127), .C2(n8292), .C3(n7442), .A(n4080), .B(N9400), 
        .ZN(n8289) );
  oan211d1 U4724 ( .C1(n8294), .C2(n8295), .B(n8296), .A(n8297), .ZN(n8292) );
  aoi31d1 U4725 ( .B1(n4088), .B2(n5036), .B3(n8299), .A(n8300), .ZN(n8294) );
  aoi311d1 U4726 ( .C1(n8301), .C2(n8302), .C3(n5943), .A(n6812), .B(n12143), 
        .ZN(n8299) );
  aoim21d1 U4727 ( .B1(images_bus[121]), .B2(n6830), .A(n7034), .ZN(n5943) );
  aon211d1 U4728 ( .C1(n4095), .C2(n8303), .B(n8304), .A(n5024), .ZN(n8301) );
  oai211d1 U4729 ( .C1(images_bus[127]), .C2(n5041), .A(n5954), .B(n8305), 
        .ZN(n8303) );
  oan211d1 U4731 ( .C1(n5948), .C2(n3996), .B(n8310), .A(n8311), .ZN(n8306) );
  aon211d1 U4732 ( .C1(n8312), .C2(images_bus[131]), .B(n8313), .A(n4004), 
        .ZN(n8310) );
  oan211d1 U4733 ( .C1(n8315), .C2(n4016), .B(n8316), .A(n5965), .ZN(n8313) );
  oan211d1 U4735 ( .C1(n5067), .C2(n8318), .B(n4015), .A(n8319), .ZN(n8316) );
  oai22d1 U4738 ( .A1(images_bus[137]), .A2(n8321), .B1(n5687), .B2(n8322), 
        .ZN(n5067) );
  aoim211d1 U4739 ( .C1(n8323), .C2(n8324), .A(n8325), .B(n8326), .ZN(n8315)
         );
  aoi31d1 U4740 ( .B1(n5970), .B2(n8327), .B3(n8324), .A(n4023), .ZN(n8326) );
  aon211d1 U4741 ( .C1(n4053), .C2(n8328), .B(n8329), .A(n4054), .ZN(n8327) );
  aon211d1 U4743 ( .C1(n4034), .C2(n8333), .B(n8334), .A(n4048), .ZN(n8331) );
  oai211d1 U4744 ( .C1(n8336), .C2(n8337), .A(n8338), .B(images_bus[153]), 
        .ZN(n8333) );
  aon211d1 U4745 ( .C1(n4039), .C2(n4959), .B(n8339), .A(n8340), .ZN(n8338) );
  aoi311d1 U4746 ( .C1(n8336), .C2(n8341), .C3(n8342), .A(n8343), .B(n8344), 
        .ZN(n8339) );
  aoi211d1 U4747 ( .C1(n3909), .C2(n8346), .A(n5112), .B(n8347), .ZN(n8342) );
  aoi22d1 U4750 ( .A1(n8350), .A2(n3917), .B1(n3916), .B2(n8353), .ZN(n8348)
         );
  oai211d1 U4751 ( .C1(n8354), .C2(n5994), .A(n8355), .B(images_bus[168]), 
        .ZN(n8353) );
  aoi211d1 U4752 ( .C1(n8356), .C2(n8357), .A(n8358), .B(n8359), .ZN(n8354) );
  ora31d1 U4753 ( .B1(n8357), .B2(n7430), .B3(n2794), .A(n8361), .Z(n8359) );
  oan211d1 U4755 ( .C1(n7429), .C2(n8363), .B(n5157), .A(n4464), .ZN(n8362) );
  oai22d1 U4756 ( .A1(n8364), .A2(n5995), .B1(n8365), .B2(n3934), .ZN(n8363)
         );
  aoi311d1 U4757 ( .C1(n3939), .C2(n5096), .C3(n8367), .A(n8368), .B(n8369), 
        .ZN(n8365) );
  oan211d1 U4759 ( .C1(n8371), .C2(n7667), .B(n3983), .A(n8373), .ZN(n8367) );
  oan211d1 U4761 ( .C1(n3961), .C2(n8375), .B(n3950), .A(n8377), .ZN(n8371) );
  oan211d1 U4762 ( .C1(n8378), .C2(n5180), .B(n5435), .A(n5773), .ZN(n8377) );
  oai22d1 U4764 ( .A1(n4958), .A2(n8380), .B1(images_bus[189]), .B2(n5772), 
        .ZN(n5184) );
  oai22d1 U4765 ( .A1(n8381), .A2(n3958), .B1(n8382), .B2(n5772), .ZN(n8379)
         );
  aoi221d1 U4767 ( .B1(n6936), .B2(n6016), .C1(n3817), .C2(n6935), .A(n8385), 
        .ZN(n8382) );
  aoi31d1 U4768 ( .B1(n8381), .B2(n5767), .B3(n8386), .A(n4431), .ZN(n8385) );
  aoi22d1 U4769 ( .A1(n3822), .A2(n8388), .B1(n8389), .B2(n3823), .ZN(n8386)
         );
  oai222d1 U4770 ( .A1(n8390), .A2(n8391), .B1(n5276), .B2(n3894), .C1(n7675), 
        .C2(n8393), .ZN(n8388) );
  aoi31d1 U4772 ( .B1(n3836), .B2(n8394), .B3(n3838), .A(n8396), .ZN(n8390) );
  oan211d1 U4773 ( .C1(n8397), .C2(n5209), .B(n3845), .A(n3837), .ZN(n8396) );
  oai22d1 U4775 ( .A1(n8401), .A2(n5214), .B1(n8402), .B2(n4409), .ZN(n8399)
         );
  oaim211d1 U4777 ( .C1(n8405), .C2(n5219), .A(n8406), .B(n8401), .ZN(n8403)
         );
  oai211d1 U4778 ( .C1(n8407), .C2(n5944), .A(n6955), .B(n3850), .ZN(n8406) );
  aoi211d1 U4779 ( .C1(n8408), .C2(n8409), .A(n4388), .B(n8410), .ZN(n8407) );
  oai211d1 U4780 ( .C1(n8411), .C2(n8412), .A(n8413), .B(n3856), .ZN(n8408) );
  aoi31d1 U4781 ( .B1(n8414), .B2(n5253), .B3(n8415), .A(n8416), .ZN(n8412) );
  aoi221d1 U4782 ( .B1(n8417), .B2(n3895), .C1(n3858), .C2(n5757), .A(n8420), 
        .ZN(n8415) );
  aoi311d1 U4783 ( .C1(n8421), .C2(n8414), .C3(n8422), .A(n8423), .B(n8424), 
        .ZN(n8420) );
  aoi22d1 U4784 ( .A1(n3863), .A2(n8426), .B1(n5257), .B2(n8082), .ZN(n8422)
         );
  oai321d1 U4785 ( .C1(n8427), .C2(n4425), .C3(n4401), .B1(n8428), .B2(n3728), 
        .A(n8429), .ZN(n8426) );
  aoi21d1 U4786 ( .B1(n3721), .B2(n8430), .A(n3619), .ZN(n8429) );
  aon211d1 U4788 ( .C1(n3807), .C2(n8431), .B(n3675), .A(n8433), .ZN(n8427) );
  oai22d1 U4790 ( .A1(images_bus[233]), .A2(n6985), .B1(n8435), .B2(n4407), 
        .ZN(n8431) );
  aoi211d1 U4791 ( .C1(n7724), .C2(n8436), .A(n8437), .B(n6989), .ZN(n8435) );
  oai21d1 U4792 ( .B1(n5182), .B2(n3806), .A(n8439), .ZN(n6989) );
  aon211d1 U4793 ( .C1(n8440), .C2(n4451), .B(n5173), .A(n3805), .ZN(n8439) );
  oai211d1 U4795 ( .C1(n8441), .C2(n8442), .A(n8443), .B(n8444), .ZN(n8436) );
  oai211d1 U4797 ( .C1(n4457), .C2(n8445), .A(images_bus[237]), .B(n5182), 
        .ZN(n6992) );
  aon211d1 U4798 ( .C1(n8446), .C2(n7003), .B(n8447), .A(n3766), .ZN(n8443) );
  aoi311d1 U4800 ( .C1(n8450), .C2(n3786), .C3(n8452), .A(n7002), .B(n3781), 
        .ZN(n8447) );
  aon211d1 U4802 ( .C1(n8453), .C2(n8454), .B(n8455), .A(n3784), .ZN(n8450) );
  aon211d1 U4803 ( .C1(n3791), .C2(n8456), .B(n5339), .A(n3678), .ZN(n8454) );
  oai31d1 U4804 ( .B1(n8458), .B2(n3577), .B3(n8455), .A(n3788), .ZN(n8456) );
  aon211d1 U4805 ( .C1(n8459), .C2(n5345), .B(n6122), .A(n4949), .ZN(n8458) );
  aoi21d1 U4806 ( .B1(n5348), .B2(n8460), .A(n8461), .ZN(n8459) );
  aoi31d1 U4808 ( .B1(images_bus[259]), .B2(n8460), .B3(n4442), .A(n8466), 
        .ZN(n8462) );
  oai211d1 U4810 ( .C1(n8469), .C2(n3515), .A(images_bus[262]), .B(n8471), 
        .ZN(n8467) );
  oan211d1 U4811 ( .C1(n8472), .C2(n7031), .B(images_bus[265]), .A(n8473), 
        .ZN(n8469) );
  aoi211d1 U4812 ( .C1(n5745), .C2(n8474), .A(n8475), .B(n3565), .ZN(n8472) );
  oai211d1 U4814 ( .C1(n8478), .C2(n4465), .A(n8479), .B(n8480), .ZN(n8474) );
  aoi211d1 U4815 ( .C1(n3538), .C2(n8481), .A(n3515), .B(n8482), .ZN(n8480) );
  aoi21d1 U4817 ( .B1(n3537), .B2(n5933), .A(n8484), .ZN(n8479) );
  aoi31d1 U4818 ( .B1(n3558), .B2(n8485), .B3(n8486), .A(n8487), .ZN(n8478) );
  oai31d1 U4819 ( .B1(n8488), .B2(n6143), .B3(n5374), .A(n8489), .ZN(n8485) );
  aon211d1 U4820 ( .C1(n3548), .C2(n8491), .B(n8492), .A(n3557), .ZN(n8488) );
  oai211d1 U4821 ( .C1(n8494), .C2(n3551), .A(n3516), .B(n3552), .ZN(n8491) );
  aoi31d1 U4824 ( .B1(n3516), .B2(n3494), .B3(n8501), .A(n8502), .ZN(n8499) );
  aoi221d1 U4825 ( .B1(n3425), .B2(n8503), .C1(n8504), .C2(n3474), .A(n8505), 
        .ZN(n8501) );
  oan211d1 U4826 ( .C1(n8506), .C2(n8507), .B(n8508), .A(n7776), .ZN(n8505) );
  aoi211d1 U4830 ( .C1(n3463), .C2(n8512), .A(n8513), .B(n3497), .ZN(n8506) );
  aon211d1 U4832 ( .C1(n8515), .C2(n3498), .B(n7783), .A(n8517), .ZN(n8513) );
  aon211d1 U4833 ( .C1(n3466), .C2(n8518), .B(n5636), .A(n3465), .ZN(n8517) );
  aoi31d1 U4835 ( .B1(n3461), .B2(n8522), .B3(n3433), .A(n7074), .ZN(n8515) );
  oai211d1 U4837 ( .C1(n8525), .C2(n8526), .A(n8527), .B(n8528), .ZN(n8522) );
  aon211d1 U4839 ( .C1(n8529), .C2(n3436), .B(n8531), .A(n3434), .ZN(n8527) );
  ora311d1 U4840 ( .C1(n8532), .C2(n3448), .C3(n8533), .A(n6184), .B(n3457), 
        .Z(n8531) );
  aon211d1 U4843 ( .C1(n7103), .C2(n8535), .B(n3442), .A(n8536), .ZN(n8533) );
  oaim211d1 U4848 ( .C1(n7110), .C2(n3446), .A(n4941), .B(n8541), .ZN(n8539)
         );
  oan211d1 U4849 ( .C1(n8542), .C2(n8543), .B(n8544), .A(n8545), .ZN(n8541) );
  oai21d1 U4850 ( .B1(n8546), .B2(n8547), .A(n3422), .ZN(n8545) );
  oan211d1 U4852 ( .C1(n8549), .C2(n3351), .B(n8551), .A(n6197), .ZN(n8543) );
  oai211d1 U4853 ( .C1(n8552), .C2(n8553), .A(n3413), .B(n3367), .ZN(n8551) );
  aoi31d1 U4854 ( .B1(n8554), .B2(n6220), .B3(n8555), .A(n6215), .ZN(n8553) );
  aoim31d1 U4855 ( .B1(n6226), .B2(n5634), .B3(n6216), .A(n8556), .ZN(n8555)
         );
  aoi211d1 U4856 ( .C1(n8557), .C2(n2795), .A(n6223), .B(n6216), .ZN(n8556) );
  oaim311d1 U4859 ( .C1(n6251), .C2(n8561), .C3(n5451), .A(n6230), .B(n6231), 
        .ZN(n8560) );
  aon211d1 U4862 ( .C1(n8566), .C2(n8567), .B(n7141), .A(n8568), .ZN(n8561) );
  aoi22d1 U4863 ( .A1(n3387), .A2(n8569), .B1(n6263), .B2(n5397), .ZN(n8566)
         );
  oai311d1 U4864 ( .C1(n8570), .C2(n8571), .C3(n8572), .A(n3392), .B(n3352), 
        .ZN(n8569) );
  aoi311d1 U4867 ( .C1(n8576), .C2(n8577), .C3(n3390), .A(n8574), .B(n4915), 
        .ZN(n8571) );
  aon211d1 U4869 ( .C1(images_bus[349]), .C2(n6281), .B(n6275), .A(n8580), 
        .ZN(n8577) );
  aon211d1 U4871 ( .C1(n4582), .C2(n8583), .B(n8584), .A(n3272), .ZN(n8582) );
  oai21d1 U4872 ( .B1(n8585), .B2(n5478), .A(n3260), .ZN(n8583) );
  aoi321d1 U4873 ( .C1(n8587), .C2(n8588), .C3(n6299), .B1(n6295), .B2(n8589), 
        .A(n8590), .ZN(n8585) );
  nd13d1 U4874 ( .A1(n8591), .A2(n8592), .A3(n6298), .ZN(n8590) );
  aor31d1 U4878 ( .B1(n8593), .B2(n4421), .B3(n8595), .A(n3282), .Z(n8594) );
  aoi22d1 U4879 ( .A1(n3286), .A2(n8597), .B1(n5487), .B2(n8598), .ZN(n8595)
         );
  aon211d1 U4880 ( .C1(n8599), .C2(n3259), .B(n5491), .A(n3259), .ZN(n8598) );
  aoi31d1 U4881 ( .B1(n8601), .B2(n8602), .B3(n3292), .A(n8604), .ZN(n8599) );
  oai211d1 U4882 ( .C1(n8605), .C2(n8606), .A(n3258), .B(n8608), .ZN(n8602) );
  oai22d1 U4885 ( .A1(n8611), .A2(n3296), .B1(n8613), .B2(n4971), .ZN(n8610)
         );
  aoi311d1 U4888 ( .C1(n3179), .C2(n8617), .C3(n8061), .A(n8618), .B(n8619), 
        .ZN(n8613) );
  nd13d1 U4890 ( .A1(n4638), .A2(n8624), .A3(n3243), .ZN(n8623) );
  oai211d1 U4891 ( .C1(n8625), .C2(n8626), .A(n8627), .B(n8628), .ZN(n8617) );
  aon211d1 U4893 ( .C1(n8632), .C2(n8633), .B(n3183), .A(n4661), .ZN(n8629) );
  aoi21d1 U4895 ( .B1(n3188), .B2(n8636), .A(n8637), .ZN(n8632) );
  oai321d1 U4896 ( .C1(n8638), .C2(n3197), .C3(n8639), .B1(n8640), .B2(n7241), 
        .A(n8641), .ZN(n8636) );
  aoi31d1 U4897 ( .B1(n8642), .B2(n5906), .B3(n3241), .A(n8643), .ZN(n8641) );
  aoi31d1 U4899 ( .B1(n3239), .B2(n8644), .B3(n8645), .A(n8646), .ZN(n8640) );
  oan211d1 U4900 ( .C1(n8647), .C2(n7247), .B(n8648), .A(n8649), .ZN(n8646) );
  oan211d1 U4901 ( .C1(n8650), .C2(n8651), .B(n8645), .A(n8652), .ZN(n8648) );
  oan211d1 U4903 ( .C1(n3233), .C2(n5806), .B(n3232), .A(n6225), .ZN(n8650) );
  oan211d1 U4904 ( .C1(n5355), .C2(n3151), .B(n8658), .A(n8659), .ZN(n8647) );
  oai22d1 U4905 ( .A1(n8660), .A2(n8661), .B1(n8658), .B2(n8662), .ZN(n8659)
         );
  oai21d1 U4906 ( .B1(n6424), .B2(n3225), .A(n8664), .ZN(n8662) );
  aoi322d1 U4907 ( .C1(n3035), .C2(n8665), .C3(n3029), .A1(n3225), .A2(n4900), 
        .B1(n3227), .B2(n8666), .ZN(n8660) );
  aon211d1 U4908 ( .C1(n3035), .C2(n3030), .B(n8668), .A(n8669), .ZN(n8666) );
  oai321d1 U4911 ( .C1(n8671), .C2(n8672), .C3(n8673), .B1(n8674), .B2(n8675), 
        .A(n8676), .ZN(n8665) );
  aoi22d1 U4912 ( .A1(n3128), .A2(n8677), .B1(n8678), .B2(n8679), .ZN(n8676)
         );
  oaim22d1 U4913 ( .A1(n8680), .A2(n8673), .B1(n8681), .B2(n8682), .ZN(n8677)
         );
  aoi31d1 U4914 ( .B1(n8683), .B2(n3052), .B3(n8684), .A(n8685), .ZN(n8674) );
  aon211d1 U4916 ( .C1(n5237), .C2(n6448), .B(n3049), .A(n8681), .ZN(n8686) );
  aoi21d1 U4918 ( .B1(n8688), .B2(images_bus[419]), .A(n6577), .ZN(n8055) );
  aoim211d1 U4919 ( .C1(n8689), .C2(n6459), .A(n6577), .B(n8690), .ZN(n8684)
         );
  aoi21d1 U4920 ( .B1(n8691), .B2(n8689), .A(n7121), .ZN(n8690) );
  oai22d1 U4921 ( .A1(images_bus[425]), .A2(n8692), .B1(n8693), .B2(n6459), 
        .ZN(n8689) );
  aoi311d1 U4922 ( .C1(n8694), .C2(n8695), .C3(n3123), .A(n8696), .B(n3067), 
        .ZN(n8693) );
  oai22d1 U4924 ( .A1(n8698), .A2(n6465), .B1(n3123), .B2(n5621), .ZN(n8696)
         );
  oan211d1 U4925 ( .C1(n8699), .C2(n7954), .B(n8700), .A(n8701), .ZN(n8698) );
  oan211d1 U4926 ( .C1(images_bus[429]), .C2(n6569), .B(n5140), .A(n3077), 
        .ZN(n8701) );
  aon211d1 U4927 ( .C1(n8703), .C2(n3121), .B(n8704), .A(n3069), .ZN(n8700) );
  aoi311d1 U4929 ( .C1(n3076), .C2(n8709), .C3(n4411), .A(n6569), .B(n8710), 
        .ZN(n8699) );
  oai22d1 U4933 ( .A1(n8712), .A2(n4408), .B1(n8714), .B2(n3119), .ZN(n8711)
         );
  aoi31d1 U4934 ( .B1(n8716), .B2(n8717), .B3(n8718), .A(n8719), .ZN(n8714) );
  oai322d1 U4936 ( .C1(n8722), .C2(n5354), .C3(n3097), .A1(n8724), .A2(n8725), 
        .B1(images_bus[440]), .B2(n3095), .ZN(n8717) );
  oan211d1 U4937 ( .C1(n6557), .C2(n8726), .B(n6554), .A(n8727), .ZN(n8724) );
  aon211d1 U4939 ( .C1(n8726), .C2(n4894), .B(n8729), .A(n8730), .ZN(n8728) );
  aoi311d1 U4940 ( .C1(n5344), .C2(n8731), .C3(n4895), .A(n8726), .B(n8733), 
        .ZN(n8729) );
  aoi311d1 U4941 ( .C1(n3017), .C2(n8734), .C3(n2927), .A(n8735), .B(n8736), 
        .ZN(n8733) );
  oan211d1 U4942 ( .C1(n2927), .C2(n8737), .B(n3105), .A(n2935), .ZN(n8735) );
  oai21d1 U4943 ( .B1(n2934), .B2(n8738), .A(n8739), .ZN(n8734) );
  aon211d1 U4944 ( .C1(n8740), .C2(n8033), .B(n8741), .A(n8738), .ZN(n8739) );
  aoi211d1 U4945 ( .C1(n8742), .C2(n8743), .A(n8744), .B(n8745), .ZN(n8741) );
  oai21d1 U4947 ( .B1(n8746), .B2(n5231), .A(n2940), .ZN(n8038) );
  aoi211d1 U4949 ( .C1(n8751), .C2(n8752), .A(n8030), .B(n8753), .ZN(n8750) );
  aoi311d1 U4950 ( .C1(n2957), .C2(n8755), .C3(N14802), .A(n8756), .B(n8752), 
        .ZN(n8753) );
  oai211d1 U4951 ( .C1(n7317), .C2(n4814), .A(n3000), .B(n8758), .ZN(n8755) );
  aoi321d1 U4952 ( .C1(n7359), .C2(n8759), .C3(n4814), .B1(n8760), .B2(n4810), 
        .A(n8761), .ZN(n8758) );
  oan211d1 U4953 ( .C1(n4405), .C2(n8763), .B(n8764), .A(n8765), .ZN(n8761) );
  aon211d1 U4954 ( .C1(n8766), .C2(n8767), .B(n8768), .A(n8763), .ZN(n8764) );
  oan211d1 U4955 ( .C1(images_bus[463]), .C2(n8769), .B(n8770), .A(n8766), 
        .ZN(n8768) );
  aoi311d1 U4957 ( .C1(images_bus[473]), .C2(n8774), .C3(n2984), .A(n8776), 
        .B(n8777), .ZN(n8773) );
  aoi211d1 U4958 ( .C1(n7356), .C2(n8778), .A(n8779), .B(n8780), .ZN(n8777) );
  oan211d1 U4959 ( .C1(images_bus[475]), .C2(n8781), .B(n8782), .A(n8783), 
        .ZN(n8780) );
  aoi31d1 U4960 ( .B1(n8782), .B2(n2984), .B3(n2976), .A(n8785), .ZN(n8779) );
  oai321d1 U4961 ( .C1(n4850), .C2(n2914), .C3(n8787), .B1(n2829), .B2(n7999), 
        .A(n8788), .ZN(n8778) );
  aoi311d1 U4962 ( .C1(n8787), .C2(n2829), .C3(n8789), .A(n8790), .B(n2817), 
        .ZN(n8788) );
  aoi211d1 U4964 ( .C1(n8793), .C2(n8794), .A(n2830), .B(n7335), .ZN(n8790) );
  oai211d1 U4967 ( .C1(n8798), .C2(n7115), .A(n8799), .B(n8800), .ZN(n8794) );
  aoi21d1 U4971 ( .B1(n4872), .B2(n7115), .A(n2865), .ZN(n8805) );
  aon211d1 U4973 ( .C1(n8807), .C2(n8808), .B(n8809), .A(n2869), .ZN(n8804) );
  oai322d1 U4974 ( .C1(n8810), .C2(images_bus[495]), .C3(n8811), .A1(n8812), 
        .A2(n8813), .B1(n4396), .B2(n2879), .ZN(n8808) );
  aoi31d1 U4976 ( .B1(n2888), .B2(n8817), .B3(n8818), .A(n8819), .ZN(n8812) );
  oai211d1 U4978 ( .C1(images_bus[504]), .C2(n2895), .A(n8822), .B(n8823), 
        .ZN(n8817) );
  oai31d1 U4979 ( .B1(n8824), .B2(n8825), .B3(n8023), .A(n2893), .ZN(n8822) );
  oai21d1 U4980 ( .B1(n4910), .B2(n4914), .A(n8826), .ZN(n8023) );
  aoi31d1 U4981 ( .B1(n4889), .B2(images_bus[504]), .B3(n4914), .A(n2898), 
        .ZN(n8825) );
  oai21d1 U4983 ( .B1(images_bus[504]), .B2(n4910), .A(n8024), .ZN(n8824) );
  aon211d1 U4985 ( .C1(n2869), .C2(n8828), .B(n4878), .A(n8829), .ZN(n7351) );
  or03d0 U4986 ( .A1(N15186), .A2(images_bus[479]), .A3(n8830), .Z(n8793) );
  oan211d1 U4987 ( .C1(n8831), .C2(n8830), .B(n8832), .A(images_bus[479]), 
        .ZN(n8789) );
  oai21d1 U4988 ( .B1(n2984), .B2(n6982), .A(n2974), .ZN(n8776) );
  or02d0 U4994 ( .A1(n8678), .A2(n6084), .Z(n8681) );
  nd13d1 U4998 ( .A1(N14162), .A2(n3037), .A3(n8680), .ZN(n8671) );
  aoi31d1 U5000 ( .B1(images_bus[407]), .B2(images_bus[406]), .B3(n8645), .A(
        n6993), .ZN(n8654) );
  oai211d1 U5003 ( .C1(n5906), .C2(n8643), .A(images_bus[400]), .B(n5518), 
        .ZN(n8639) );
  aoi31d1 U5008 ( .B1(n8619), .B2(images_bus[390]), .B3(images_bus[391]), .A(
        n7127), .ZN(n8628) );
  or02d0 U5010 ( .A1(n8834), .A2(n4970), .Z(n8618) );
  aon211d1 U5012 ( .C1(n3237), .C2(images_bus[403]), .B(n8836), .A(n3205), 
        .ZN(n8638) );
  oai22d1 U5015 ( .A1(n8838), .A2(n7197), .B1(n8839), .B2(n8616), .ZN(n4631)
         );
  oai211d1 U5016 ( .C1(n8840), .C2(n8616), .A(n8608), .B(n7198), .ZN(n8609) );
  aoi211d1 U5017 ( .C1(n8834), .C2(n8062), .A(n8064), .B(n8063), .ZN(n8840) );
  oai21d1 U5018 ( .B1(n8841), .B2(n8842), .A(n8843), .ZN(n8064) );
  oai21d1 U5019 ( .B1(n8844), .B2(n8842), .A(n8845), .ZN(n8062) );
  aon211d1 U5035 ( .C1(images_bus[363]), .C2(n4601), .B(n7381), .A(n7382), 
        .ZN(n8587) );
  aoim31d1 U5038 ( .B1(n8568), .B2(n12157), .B3(n5825), .A(n6998), .ZN(n8567)
         );
  aoi321d1 U5041 ( .C1(n6232), .C2(n5927), .C3(n8848), .B1(n8564), .B2(n8846), 
        .A(n8849), .ZN(n8557) );
  nd13d1 U5042 ( .A1(n8849), .A2(n6602), .A3(images_bus[335]), .ZN(n8846) );
  aoi21d1 U5047 ( .B1(n5633), .B2(n3410), .A(n8851), .ZN(n6220) );
  aoi21d1 U5050 ( .B1(images_bus[327]), .B2(n8552), .A(n7136), .ZN(n8554) );
  aoi31d1 U5058 ( .B1(n8529), .B2(images_bus[311]), .B3(n4308), .A(n7006), 
        .ZN(n8536) );
  oai21d1 U5059 ( .B1(n3345), .B2(n8854), .A(n4941), .ZN(n7110) );
  aoi31d1 U5066 ( .B1(n5735), .B2(images_bus[295]), .B3(n8504), .A(n7150), 
        .ZN(n8508) );
  oai31d1 U5071 ( .B1(n8489), .B2(n6242), .B3(n5834), .A(images_bus[280]), 
        .ZN(n8492) );
  aoim21d1 U5073 ( .B1(n5933), .B2(n8481), .A(n5740), .ZN(n8487) );
  aoi21d1 U5075 ( .B1(n8460), .B2(n4681), .A(n7152), .ZN(n8483) );
  oai21d1 U5088 ( .B1(n4949), .B2(n7013), .A(images_bus[251]), .ZN(n5342) );
  aoi31d1 U5093 ( .B1(n8859), .B2(n5748), .B3(n4692), .A(n12118), .ZN(n8434)
         );
  aoi21d1 U5098 ( .B1(n4951), .B2(n3857), .A(n3860), .ZN(n5253) );
  aoi21d1 U5100 ( .B1(n8862), .B2(n8411), .A(n7019), .ZN(n8414) );
  oai211d1 U5102 ( .C1(n5944), .C2(n8405), .A(images_bus[208]), .B(n5550), 
        .ZN(n8409) );
  nd13d1 U5103 ( .A1(n8394), .A2(n8864), .A3(n8401), .ZN(n8405) );
  oai31d1 U5104 ( .B1(n8393), .B2(n6390), .B3(n6038), .A(images_bus[200]), 
        .ZN(n8394) );
  aoi21d1 U5106 ( .B1(n5767), .B2(n8381), .A(n5766), .ZN(n8389) );
  oaim21d1 U5108 ( .B1(n8865), .B2(n8369), .A(images_bus[184]), .ZN(n8375) );
  aor31d1 U5119 ( .B1(n4320), .B2(n8328), .B3(n5570), .A(n7023), .Z(n8334) );
  oai21d1 U5124 ( .B1(images_bus[141]), .B2(n5074), .A(images_bus[139]), .ZN(
        n8325) );
  oai21d1 U5126 ( .B1(n6647), .B2(n3996), .A(images_bus[136]), .ZN(n8318) );
  aoi21d1 U5130 ( .B1(images_bus[127]), .B2(n8308), .A(n5053), .ZN(n8312) );
  aon211d1 U5139 ( .C1(n4097), .C2(n8875), .B(n4965), .A(n8876), .ZN(n8874) );
  aoi211d1 U5153 ( .C1(n7447), .C2(n4167), .A(n8881), .B(n5456), .ZN(n5868) );
  aoi31d1 U5155 ( .B1(n4323), .B2(n5852), .B3(n8882), .A(n7042), .ZN(n8264) );
  aoi311d1 U5156 ( .C1(images_bus[79]), .C2(n4510), .C3(n4219), .A(n6662), .B(
        n7104), .ZN(n8882) );
  oai21d1 U5161 ( .B1(n6748), .B2(n8243), .A(n5697), .ZN(n8246) );
  aoi21d1 U5164 ( .B1(images_bus[63]), .B2(n8233), .A(n5807), .ZN(n8238) );
  nd13d1 U5167 ( .A1(n8207), .A2(n4330), .A3(images_bus[55]), .ZN(n8220) );
  oai31d1 U5172 ( .B1(n8887), .B2(n6070), .B3(n6694), .A(images_bus[40]), .ZN(
        n8187) );
  oai21d1 U5179 ( .B1(n7481), .B2(n8157), .A(images_bus[24]), .ZN(n8162) );
  oai21d1 U5180 ( .B1(n5964), .B2(n4523), .A(n7477), .ZN(n8157) );
  aoi21d1 U5187 ( .B1(images_bus[4]), .B2(n8890), .A(n7461), .ZN(N26360) );
  aon211d1 U5188 ( .C1(n4858), .C2(n8892), .B(n8893), .A(n8894), .ZN(n8890) );
  aon211d1 U5189 ( .C1(n8895), .C2(images_bus[6]), .B(n7586), .A(n8897), .ZN(
        n8892) );
  aoi22d1 U5191 ( .A1(n4766), .A2(n8899), .B1(n8900), .B2(n8901), .ZN(n8895)
         );
  oai22d1 U5192 ( .A1(n4866), .A2(n8903), .B1(n8904), .B2(n8144), .ZN(n8899)
         );
  aoi31d1 U5194 ( .B1(n4819), .B2(n8906), .B3(n4816), .A(n8907), .ZN(n8904) );
  oai311d1 U5195 ( .C1(n7462), .C2(n8908), .C3(n8909), .A(n8910), .B(
        images_bus[13]), .ZN(n8906) );
  aon211d1 U5196 ( .C1(n4604), .C2(n4530), .B(n6355), .A(n4628), .ZN(n8910) );
  aoi321d1 U5197 ( .C1(n4392), .C2(n8914), .C3(n4552), .B1(n4561), .B2(n4524), 
        .A(n8918), .ZN(n8908) );
  oai22d1 U5198 ( .A1(images_bus[21]), .A2(n8919), .B1(n8920), .B2(n7473), 
        .ZN(n8918) );
  oai211d1 U5201 ( .C1(images_bus[22]), .C2(n8922), .A(n8921), .B(n8923), .ZN(
        n8914) );
  aoi22d1 U5202 ( .A1(n8924), .A2(n4373), .B1(n4357), .B2(n8926), .ZN(n8923)
         );
  oan211d1 U5203 ( .C1(n8927), .C2(n8125), .B(n8928), .A(n6679), .ZN(n8924) );
  aoi31d1 U5205 ( .B1(n7487), .B2(n8926), .B3(images_bus[24]), .A(n7494), .ZN(
        n8928) );
  oai21d1 U5208 ( .B1(images_bus[31]), .B2(n6671), .A(n8176), .ZN(n8123) );
  aoi31d1 U5209 ( .B1(n2792), .B2(n8126), .B3(n8933), .A(n6671), .ZN(n8931) );
  oan211d1 U5211 ( .C1(n8936), .C2(n8937), .B(n8938), .A(n7496), .ZN(n8935) );
  aon211d1 U5212 ( .C1(n4276), .C2(n8940), .B(n4754), .A(n4233), .ZN(n8938) );
  oai211d1 U5213 ( .C1(n8942), .C2(n8943), .A(images_bus[37]), .B(n8936), .ZN(
        n8940) );
  aoi211d1 U5214 ( .C1(n5788), .C2(n8944), .A(n8945), .B(n4246), .ZN(n8942) );
  oai322d1 U5215 ( .C1(n5704), .C2(n8946), .C3(n7183), .A1(n8947), .A2(n6710), 
        .B1(n6711), .B2(n8948), .ZN(n8944) );
  oan211d1 U5216 ( .C1(n8949), .C2(n8950), .B(n8197), .A(n8951), .ZN(n8947) );
  aoi31d1 U5217 ( .B1(n4285), .B2(n8953), .B3(n6714), .A(n8954), .ZN(n8949) );
  aoi21d1 U5220 ( .B1(n8958), .B2(n8959), .A(n8204), .ZN(n8955) );
  oai211d1 U5222 ( .C1(n8963), .C2(n8964), .A(n8965), .B(n4284), .ZN(n8962) );
  aoi211d1 U5223 ( .C1(n8967), .C2(n8968), .A(n8969), .B(n8970), .ZN(n8963) );
  oai321d1 U5224 ( .C1(n8971), .C2(n8972), .C3(n8215), .B1(n8973), .B2(n8974), 
        .A(n4331), .ZN(n8969) );
  aoi31d1 U5225 ( .B1(images_bus[56]), .B2(n4283), .B3(images_bus[57]), .A(
        n8976), .ZN(n8972) );
  oan211d1 U5226 ( .C1(n8973), .C2(n8977), .B(n8978), .A(n8979), .ZN(n8976) );
  oai211d1 U5227 ( .C1(n8980), .C2(n4282), .A(n4266), .B(n8983), .ZN(n8978) );
  oan211d1 U5229 ( .C1(n8985), .C2(n8986), .B(n8984), .A(n4267), .ZN(n8980) );
  oan211d1 U5231 ( .C1(n8989), .C2(n8990), .B(n8991), .A(n6733), .ZN(n8985) );
  oai21d1 U5232 ( .B1(n8884), .B2(n8992), .A(images_bus[61]), .ZN(n6733) );
  oai22d1 U5233 ( .A1(n8235), .A2(n8993), .B1(n8994), .B2(n8995), .ZN(n8990)
         );
  aoi31d1 U5234 ( .B1(n4187), .B2(n8996), .B3(n4188), .A(n8998), .ZN(n8994) );
  oan211d1 U5235 ( .C1(n8999), .C2(n9000), .B(n4184), .A(n4185), .ZN(n8998) );
  oai21d1 U5239 ( .B1(images_bus[71]), .B2(n9004), .A(n9005), .ZN(n9003) );
  aon211d1 U5240 ( .C1(n4149), .C2(n9006), .B(n9007), .A(n9008), .ZN(n9005) );
  oai222d1 U5241 ( .A1(n9009), .A2(n5039), .B1(n9010), .B2(n9011), .C1(n9012), 
        .C2(n9013), .ZN(n9006) );
  oan211d1 U5242 ( .C1(n9014), .C2(n8251), .B(n4180), .A(n9015), .ZN(n9009) );
  aoi31d1 U5243 ( .B1(n4142), .B2(n5840), .B3(n9017), .A(n4155), .ZN(n9014) );
  aoi22d1 U5244 ( .A1(n9018), .A2(n9019), .B1(n9020), .B2(n5023), .ZN(n9017)
         );
  oaim22d1 U5245 ( .A1(n8259), .A2(n9021), .B1(n5023), .B2(n9022), .ZN(n9019)
         );
  oan211d1 U5246 ( .C1(n6768), .C2(images_bus[85]), .B(n9023), .A(n5853), .ZN(
        n9022) );
  aon211d1 U5249 ( .C1(n4163), .C2(n9024), .B(n4326), .A(n7548), .ZN(n9021) );
  aoi21d1 U5251 ( .B1(n4172), .B2(n9027), .A(n9028), .ZN(n9025) );
  aoi321d1 U5252 ( .C1(images_bus[93]), .C2(n9029), .C3(n4141), .B1(n4141), 
        .B2(n5027), .A(n5037), .ZN(n9028) );
  oai211d1 U5254 ( .C1(n9032), .C2(n5879), .A(n9033), .B(n4118), .ZN(n9029) );
  oai211d1 U5255 ( .C1(n5882), .C2(n9035), .A(n9036), .B(n9037), .ZN(n9033) );
  aon211d1 U5256 ( .C1(n9038), .C2(n4063), .B(n9040), .A(n4115), .ZN(n9036) );
  oan211d1 U5258 ( .C1(n9044), .C2(n6786), .B(images_bus[101]), .A(n5019), 
        .ZN(n9038) );
  aoi321d1 U5259 ( .C1(n4111), .C2(n9046), .C3(n4068), .B1(n6787), .B2(n9048), 
        .A(n9049), .ZN(n9044) );
  oai21d1 U5260 ( .B1(n9042), .B2(n9050), .A(n4070), .ZN(n9049) );
  oai21d1 U5262 ( .B1(images_bus[102]), .B2(n9050), .A(images_bus[101]), .ZN(
        n6789) );
  oaim31d1 U5263 ( .B1(images_bus[105]), .B2(n9048), .B3(images_bus[104]), .A(
        n9052), .ZN(n9046) );
  oai211d1 U5264 ( .C1(n9053), .C2(n9054), .A(n5909), .B(n4073), .ZN(n9052) );
  aoi31d1 U5265 ( .B1(n4137), .B2(n6800), .B3(n9057), .A(n8290), .ZN(n9053) );
  aoi31d1 U5266 ( .B1(n4077), .B2(n4081), .B3(n9060), .A(n4076), .ZN(n9057) );
  aoim21d1 U5268 ( .B1(n9063), .B2(n4085), .A(n9065), .ZN(n9060) );
  oan211d1 U5271 ( .C1(n9070), .C2(n5940), .B(images_bus[117]), .A(n5935), 
        .ZN(n9067) );
  aoi321d1 U5273 ( .C1(n9073), .C2(n4091), .C3(n9075), .B1(n9076), .B2(n9077), 
        .A(n5936), .ZN(n9070) );
  aoi21d1 U5274 ( .B1(n9078), .B2(n9079), .A(n6835), .ZN(n9075) );
  oai211d1 U5276 ( .C1(n3991), .C2(n5041), .A(images_bus[125]), .B(n9083), 
        .ZN(n9082) );
  aoi221d1 U5277 ( .B1(n3999), .B2(n4136), .C1(n3999), .C2(n6649), .A(n9085), 
        .ZN(n9083) );
  oan211d1 U5278 ( .C1(n5948), .C2(n9086), .B(n9087), .A(n3998), .ZN(n9085) );
  oai211d1 U5280 ( .C1(n5056), .C2(n9088), .A(n4056), .B(n4391), .ZN(n9087) );
  oai21d1 U5281 ( .B1(n5281), .B2(n9086), .A(n9090), .ZN(n9088) );
  aon211d1 U5282 ( .C1(n4008), .C2(n9092), .B(n9093), .A(n4014), .ZN(n9090) );
  aoi31d1 U5283 ( .B1(n3990), .B2(images_bus[134]), .B3(n9096), .A(n5007), 
        .ZN(n9093) );
  aoi22d1 U5284 ( .A1(n9097), .A2(n7614), .B1(n9098), .B2(n9099), .ZN(n9096)
         );
  oan211d1 U5285 ( .C1(n9100), .C2(n9101), .B(n9102), .A(n8323), .ZN(n9097) );
  aon211d1 U5286 ( .C1(n4025), .C2(n9103), .B(n4491), .A(n9104), .ZN(n9101) );
  aon211d1 U5287 ( .C1(n9105), .C2(images_bus[143]), .B(n5076), .A(n5077), 
        .ZN(n9103) );
  aoi22d1 U5288 ( .A1(n4051), .A2(n9107), .B1(n9108), .B2(n4027), .ZN(n9105)
         );
  oaim31d1 U5289 ( .B1(n4027), .B2(n12144), .B3(n5088), .A(n9110), .ZN(n9107)
         );
  aon211d1 U5290 ( .C1(n4048), .C2(n9111), .B(n4319), .A(n6854), .ZN(n9110) );
  oai321d1 U5291 ( .C1(n9112), .C2(n8343), .C3(n7437), .B1(n9113), .B2(n4389), 
        .A(n9114), .ZN(n9111) );
  aoi21d1 U5293 ( .B1(n8096), .B2(n4047), .A(n4319), .ZN(n5092) );
  aon211d1 U5294 ( .C1(n4044), .C2(n9118), .B(n9119), .A(n8340), .ZN(n9112) );
  oai321d1 U5295 ( .C1(n4418), .C2(n9120), .C3(n6874), .B1(n8869), .B2(n5115), 
        .A(n9121), .ZN(n9118) );
  aoi21d1 U5298 ( .B1(n7645), .B2(n7647), .A(n9122), .ZN(n8341) );
  aoi221d1 U5299 ( .B1(n6883), .B2(n9123), .C1(n3917), .C2(n4703), .A(n9124), 
        .ZN(n9120) );
  aoi311d1 U5300 ( .C1(n3981), .C2(n4719), .C3(n9126), .A(n6880), .B(n7652), 
        .ZN(n9124) );
  aoi22d1 U5301 ( .A1(n8867), .A2(n9127), .B1(n3922), .B2(n9128), .ZN(n9126)
         );
  oai22d1 U5302 ( .A1(n9129), .A2(n4422), .B1(n9130), .B2(n5144), .ZN(n9127)
         );
  aoi322d1 U5303 ( .C1(images_bus[169]), .C2(n9128), .C3(images_bus[168]), 
        .A1(n7654), .A2(n9131), .B1(n3931), .B2(n9132), .ZN(n9130) );
  oai321d1 U5306 ( .C1(n3934), .C2(n9133), .C3(n8373), .B1(n3978), .B2(n5995), 
        .A(n4470), .ZN(n9131) );
  aoi221d1 U5308 ( .B1(n3939), .B2(n9137), .C1(n5170), .C2(n9138), .A(n5172), 
        .ZN(n9133) );
  oai222d1 U5310 ( .A1(n9140), .A2(n5773), .B1(n3979), .B2(n3946), .C1(n4317), 
        .C2(n7428), .ZN(n9138) );
  aoi211d1 U5314 ( .C1(n3957), .C2(n9145), .A(n9146), .B(n9147), .ZN(n9140) );
  oai21d1 U5315 ( .B1(n9148), .B2(n6009), .A(n9149), .ZN(n9146) );
  aoi31d1 U5318 ( .B1(n3828), .B2(n9150), .B3(n3823), .A(n9151), .ZN(n9148) );
  oai22d1 U5319 ( .A1(n9152), .A2(n9153), .B1(n9154), .B2(n5198), .ZN(n9150)
         );
  aon211d1 U5321 ( .C1(n5201), .C2(n9156), .B(n12170), .A(n3835), .ZN(n9152)
         );
  oai211d1 U5322 ( .C1(n3892), .C2(n5206), .A(n9154), .B(n9158), .ZN(n9156) );
  aoi221d1 U5323 ( .B1(n5211), .B2(n9159), .C1(n3880), .C2(n6390), .A(n12170), 
        .ZN(n9158) );
  oai322d1 U5324 ( .C1(n5669), .C2(n3892), .C3(n7155), .A1(n9160), .A2(n9161), 
        .B1(n3893), .B2(n4409), .ZN(n9159) );
  aon211d1 U5328 ( .C1(n3877), .C2(n9166), .B(n4459), .A(n9167), .ZN(n9160) );
  oai321d1 U5329 ( .C1(n5230), .C2(n9168), .C3(n8410), .B1(n9169), .B2(n5227), 
        .A(n9170), .ZN(n9166) );
  aoi31d1 U5331 ( .B1(n3873), .B2(n9172), .B3(n8413), .A(n9173), .ZN(n9168) );
  oai211d1 U5332 ( .C1(n9174), .C2(n7417), .A(n9175), .B(n9176), .ZN(n9172) );
  aoi211d1 U5333 ( .C1(n5240), .C2(n7704), .A(n9177), .B(n4314), .ZN(n9174) );
  aor22d1 U5334 ( .A1(n9178), .A2(n3868), .B1(n9180), .B2(n4412), .Z(n9177) );
  aor31d1 U5335 ( .B1(n5257), .B2(n9181), .B3(n3865), .A(n9183), .Z(n9180) );
  aoi211d1 U5337 ( .C1(n3721), .C2(n7711), .A(n3619), .B(n9186), .ZN(n9184) );
  oan211d1 U5338 ( .C1(n9187), .C2(n3730), .B(images_bus[223]), .A(n3728), 
        .ZN(n9186) );
  aoi22d1 U5340 ( .A1(n3744), .A2(n9190), .B1(n9191), .B2(n3736), .ZN(n9187)
         );
  oai321d1 U5341 ( .C1(n5287), .C2(n9193), .C3(n5286), .B1(images_bus[229]), 
        .B2(n9194), .A(n9195), .ZN(n9190) );
  oai311d1 U5342 ( .C1(n9196), .C2(n9197), .C3(n3719), .A(n9199), .B(n3738), 
        .ZN(n9195) );
  oai21d1 U5343 ( .B1(n9201), .B2(n9202), .A(n9203), .ZN(n9196) );
  oan211d1 U5345 ( .C1(n9207), .C2(n3806), .B(n3712), .A(n9209), .ZN(n9206) );
  aon211d1 U5347 ( .C1(n9213), .C2(n5303), .B(n5305), .A(n9214), .ZN(n9210) );
  aon211d1 U5348 ( .C1(n3801), .C2(n9215), .B(n5308), .A(n5309), .ZN(n9213) );
  oai211d1 U5349 ( .C1(n5317), .C2(n9216), .A(n9217), .B(images_bus[239]), 
        .ZN(n9215) );
  oai211d1 U5350 ( .C1(n9218), .C2(n9219), .A(n3777), .B(n6999), .ZN(n9217) );
  oan211d1 U5352 ( .C1(n9220), .C2(n9221), .B(images_bus[245]), .A(n9222), 
        .ZN(n9218) );
  aoi211d1 U5353 ( .C1(n9223), .C2(n9224), .A(n9219), .B(n4313), .ZN(n9220) );
  oai321d1 U5354 ( .C1(n3781), .C2(n9225), .C3(n5334), .B1(n9226), .B2(n9227), 
        .A(n8857), .ZN(n9224) );
  aoi31d1 U5355 ( .B1(n5337), .B2(n3790), .B3(n9229), .A(n9230), .ZN(n9225) );
  oan211d1 U5358 ( .C1(n9231), .C2(n7015), .B(n9232), .A(n5339), .ZN(n9229) );
  aoi311d1 U5359 ( .C1(n3789), .C2(n9233), .C3(n3575), .A(n3715), .B(n7020), 
        .ZN(n9231) );
  aoi22d1 U5363 ( .A1(n7027), .A2(n9237), .B1(n5348), .B2(n9238), .ZN(n9236)
         );
  oai211d1 U5364 ( .C1(images_bus[261]), .C2(n9239), .A(n9240), .B(n9241), 
        .ZN(n9237) );
  aoi221d1 U5366 ( .B1(n8471), .B2(n9244), .C1(n5744), .C2(n9245), .A(n6388), 
        .ZN(n9242) );
  oai211d1 U5367 ( .C1(n9246), .C2(n9247), .A(n9248), .B(n9249), .ZN(n9245) );
  aoi211d1 U5368 ( .C1(n9250), .C2(n7406), .A(n9251), .B(n9252), .ZN(n9249) );
  aoi211d1 U5370 ( .C1(n9255), .C2(n9256), .A(n9257), .B(n6533), .ZN(n9253) );
  oai22d1 U5371 ( .A1(n4312), .A2(n9259), .B1(n9260), .B2(n9261), .ZN(n9257)
         );
  aoi321d1 U5372 ( .C1(n3547), .C2(n6154), .C3(n9263), .B1(n9264), .B2(n3549), 
        .A(n5834), .ZN(n9260) );
  oan211d1 U5373 ( .C1(n6165), .C2(n9266), .B(n9267), .A(n9268), .ZN(n9263) );
  aon211d1 U5374 ( .C1(n9269), .C2(n3477), .B(n3478), .A(n3556), .ZN(n9266) );
  aoi22d1 U5375 ( .A1(n3490), .A2(n9271), .B1(n9272), .B2(n9273), .ZN(n9269)
         );
  oai211d1 U5376 ( .C1(n3493), .C2(n9275), .A(n9276), .B(n9277), .ZN(n9271) );
  aoi211d1 U5377 ( .C1(n9278), .C2(n9279), .A(n8510), .B(n12122), .ZN(n9275)
         );
  oai211d1 U5378 ( .C1(n9280), .C2(n9281), .A(n9282), .B(n3473), .ZN(n9278) );
  aon211d1 U5379 ( .C1(n9283), .C2(n3426), .B(n6169), .A(n9285), .ZN(n9282) );
  oai211d1 U5380 ( .C1(n6169), .C2(n3426), .A(images_bus[293]), .B(n9283), 
        .ZN(n9281) );
  oai322d1 U5382 ( .C1(n4495), .C2(n9286), .C3(n5396), .A1(n9287), .A2(n5392), 
        .B1(n3491), .B2(n9289), .ZN(n9280) );
  aoi31d1 U5384 ( .B1(images_bus[296]), .B2(n9290), .B3(images_bus[297]), .A(
        n9291), .ZN(n9286) );
  aoi211d1 U5385 ( .C1(n9292), .C2(n9293), .A(n9294), .B(n5402), .ZN(n9291) );
  oai31d1 U5386 ( .B1(n9295), .B2(n8523), .B3(n9296), .A(n3461), .ZN(n9293) );
  aoi31d1 U5387 ( .B1(n9292), .B2(images_bus[303]), .B3(n9297), .A(n5404), 
        .ZN(n9296) );
  aoi211d1 U5388 ( .C1(n9298), .C2(n3435), .A(n9299), .B(n9300), .ZN(n9297) );
  aoi311d1 U5389 ( .C1(n9301), .C2(n7094), .C3(n9302), .A(n9303), .B(n7090), 
        .ZN(n9300) );
  oaim31d1 U5391 ( .B1(n9302), .B2(images_bus[309]), .B3(n9305), .A(n7091), 
        .ZN(n9301) );
  aoi31d1 U5393 ( .B1(n3449), .B2(n9306), .B3(n7100), .A(n9307), .ZN(n9305) );
  oan211d1 U5394 ( .C1(n3492), .C2(n9309), .B(n4308), .A(n9310), .ZN(n9307) );
  aon211d1 U5397 ( .C1(n9313), .C2(n9314), .B(n9315), .A(n9316), .ZN(n9306) );
  oai211d1 U5399 ( .C1(n6188), .C2(n9317), .A(n9318), .B(n6194), .ZN(n9313) );
  oaim21d1 U5400 ( .B1(n9317), .B2(n9319), .A(n9320), .ZN(n9318) );
  oai321d1 U5401 ( .C1(n8854), .C2(n9321), .C3(n5418), .B1(n3340), .B2(n8547), 
        .A(n9323), .ZN(n9317) );
  aoi31d1 U5402 ( .B1(n3364), .B2(n9325), .B3(n8544), .A(n7812), .ZN(n9323) );
  oai311d1 U5404 ( .C1(n7817), .C2(n9326), .C3(n3412), .A(n9328), .B(n9329), 
        .ZN(n9325) );
  aon211d1 U5405 ( .C1(n3416), .C2(n4663), .B(n9331), .A(n3367), .ZN(n9329) );
  aoi211d1 U5406 ( .C1(n3414), .C2(n9332), .A(n9331), .B(n4663), .ZN(n9326) );
  oai321d1 U5407 ( .C1(n9333), .C2(n9334), .C3(n6215), .B1(n3341), .B2(n9336), 
        .A(n9337), .ZN(n9332) );
  aoi321d1 U5408 ( .C1(n3409), .C2(n9338), .C3(n3405), .B1(n7818), .B2(n9339), 
        .A(n9340), .ZN(n9334) );
  oai221d1 U5411 ( .B1(images_bus[333]), .B2(n9342), .C1(n9343), .C2(n3403), 
        .A(n3344), .ZN(n9339) );
  aoi221d1 U5414 ( .B1(n6232), .B2(n9347), .C1(n3375), .C2(n9348), .A(n9349), 
        .ZN(n9343) );
  oai222d1 U5415 ( .A1(n9350), .A2(n3378), .B1(n8850), .B2(n9352), .C1(n3343), 
        .C2(n9354), .ZN(n9348) );
  aoi22d1 U5416 ( .A1(n9355), .A2(n9356), .B1(n7135), .B2(n9357), .ZN(n9350)
         );
  oai221d1 U5417 ( .B1(n3343), .B2(n5455), .C1(n9358), .C2(n6258), .A(
        images_bus[341]), .ZN(n9357) );
  aoi221d1 U5418 ( .B1(n9359), .B2(n3394), .C1(n3397), .C2(n3342), .A(n9361), 
        .ZN(n9358) );
  oan211d1 U5419 ( .C1(n9362), .C2(n9363), .B(n9364), .A(n5462), .ZN(n9359) );
  aoi311d1 U5421 ( .C1(n7850), .C2(n3271), .C3(n9365), .A(n9366), .B(n9367), 
        .ZN(n9362) );
  oan211d1 U5422 ( .C1(n3261), .C2(n4579), .B(n3251), .A(n9369), .ZN(n9367) );
  oai21d1 U5424 ( .B1(n9371), .B2(n7841), .A(n9372), .ZN(n9366) );
  aoim21d1 U5425 ( .B1(n5463), .B2(n3391), .A(n9373), .ZN(n7841) );
  aoi21d1 U5426 ( .B1(n9374), .B2(n8581), .A(n9369), .ZN(n9373) );
  oan211d1 U5427 ( .C1(n9375), .C2(n9376), .B(n9377), .A(n9369), .ZN(n9365) );
  aoi321d1 U5428 ( .C1(n6292), .C2(n3321), .C3(n9378), .B1(n6292), .B2(n9379), 
        .A(n9380), .ZN(n9375) );
  oai21d1 U5429 ( .B1(n9381), .B2(n4586), .A(n9377), .ZN(n9380) );
  aoi31d1 U5430 ( .B1(n9381), .B2(n4656), .B3(n9382), .A(n9379), .ZN(n9378) );
  aoi321d1 U5431 ( .C1(n6314), .C2(n5480), .C3(n9383), .B1(n3319), .B2(n9385), 
        .A(n6301), .ZN(n9382) );
  aoi311d1 U5432 ( .C1(n9386), .C2(n3286), .C3(n9387), .A(n9388), .B(n9389), 
        .ZN(n9383) );
  aoi21d1 U5433 ( .B1(n3283), .B2(n9390), .A(n9391), .ZN(n9389) );
  aon211d1 U5434 ( .C1(n9386), .C2(n4421), .B(n3282), .A(n6311), .ZN(n9390) );
  oan211d1 U5438 ( .C1(n9395), .C2(n9396), .B(n3292), .A(n9397), .ZN(n9393) );
  oai21d1 U5440 ( .B1(images_bus[373]), .B2(n9398), .A(n9399), .ZN(n9396) );
  oai222d1 U5441 ( .A1(n9400), .A2(n9401), .B1(n4305), .B2(n9402), .C1(n3262), 
        .C2(n9404), .ZN(n9395) );
  aoim211d1 U5443 ( .C1(n6593), .C2(n8841), .A(n9406), .B(n9407), .ZN(n9400)
         );
  aoi31d1 U5444 ( .B1(n3146), .B2(n9408), .B3(n3263), .A(n9410), .ZN(n9407) );
  oai211d1 U5446 ( .C1(n3150), .C2(n9412), .A(n3250), .B(n3248), .ZN(n9408) );
  oan211d1 U5447 ( .C1(n9415), .C2(n8621), .B(n9416), .A(n3246), .ZN(n9412) );
  aoi321d1 U5448 ( .C1(n3178), .C2(n3177), .C3(n9420), .B1(n9421), .B2(n9422), 
        .A(n9423), .ZN(n9415) );
  oan211d1 U5449 ( .C1(n5242), .C2(n9416), .B(n6600), .A(n8620), .ZN(n9423) );
  oan211d1 U5450 ( .C1(n9424), .C2(n6377), .B(images_bus[390]), .A(n8620), 
        .ZN(n9420) );
  aoi31d1 U5451 ( .B1(n9425), .B2(n9426), .B3(n3243), .A(n5982), .ZN(n9424) );
  oai31d1 U5452 ( .B1(n9427), .B2(n6379), .B3(n9428), .A(images_bus[391]), 
        .ZN(n9426) );
  aon211d1 U5453 ( .C1(n9429), .C2(n9430), .B(n6558), .A(n9431), .ZN(n9427) );
  or02d0 U5454 ( .A1(n9430), .A2(n6391), .Z(n9431) );
  oai211d1 U5455 ( .C1(n4964), .C2(n6391), .A(n8635), .B(n9432), .ZN(n9430) );
  aon211d1 U5456 ( .C1(n8642), .C2(n5906), .B(n9433), .A(n6386), .ZN(n9432) );
  oaim211d1 U5459 ( .C1(n9435), .C2(n6401), .A(n3199), .B(n3195), .ZN(n9434)
         );
  aoi21d1 U5460 ( .B1(n9438), .B2(images_bus[403]), .A(n8836), .ZN(n6401) );
  oai321d1 U5462 ( .C1(n6409), .C2(images_bus[405]), .C3(n3235), .B1(
        images_bus[404]), .B2(n3207), .A(n9441), .ZN(n9440) );
  aon211d1 U5463 ( .C1(n3211), .C2(n9442), .B(n9443), .A(n3207), .ZN(n9441) );
  oan211d1 U5464 ( .C1(n9444), .C2(n9445), .B(n9446), .A(n7247), .ZN(n9443) );
  oai21d1 U5467 ( .B1(n3227), .B2(n4900), .A(n3222), .ZN(n7374) );
  aoi221d1 U5469 ( .B1(n9449), .B2(n12150), .C1(n3032), .C2(n9451), .A(n3018), 
        .ZN(n9444) );
  oai222d1 U5472 ( .A1(n8675), .A2(n9454), .B1(n8679), .B2(n9455), .C1(n5706), 
        .C2(n3128), .ZN(n9451) );
  aon211d1 U5473 ( .C1(images_bus[416]), .C2(n6578), .B(n7919), .A(n6084), 
        .ZN(n9455) );
  aon211d1 U5474 ( .C1(n4715), .C2(n9456), .B(n9457), .A(n3050), .ZN(n9454) );
  oan211d1 U5475 ( .C1(n9459), .C2(n3047), .B(n4720), .A(n6599), .ZN(n9457) );
  oai22d1 U5476 ( .A1(images_bus[421]), .A2(n9459), .B1(n9461), .B2(n9462), 
        .ZN(n9456) );
  aon211d1 U5477 ( .C1(n7948), .C2(n4953), .B(n9463), .A(n9459), .ZN(n9462) );
  oan211d1 U5478 ( .C1(images_bus[423]), .C2(n9464), .B(n9465), .A(n7948), 
        .ZN(n9463) );
  oai211d1 U5479 ( .C1(n9466), .C2(n9467), .A(n7939), .B(n3058), .ZN(n9465) );
  oan211d1 U5482 ( .C1(n6556), .C2(n5589), .B(n9470), .A(n9471), .ZN(n9466) );
  oai21d1 U5483 ( .B1(n9472), .B2(n9473), .A(n3064), .ZN(n9470) );
  aon211d1 U5484 ( .C1(n3073), .C2(n5703), .B(n6556), .A(n9474), .ZN(n9473) );
  aon211d1 U5485 ( .C1(n6468), .C2(n6568), .B(n9475), .A(n3072), .ZN(n9474) );
  aoi311d1 U5488 ( .C1(n3103), .C2(n9481), .C3(n3100), .A(n9482), .B(n9483), 
        .ZN(n9479) );
  aoi311d1 U5489 ( .C1(n9484), .C2(n9485), .C3(n3110), .A(n6487), .B(
        images_bus[439]), .ZN(n9483) );
  oan211d1 U5491 ( .C1(n3102), .C2(n4894), .B(n3106), .A(n6990), .ZN(n9487) );
  oai21d1 U5494 ( .B1(n6559), .B2(n8722), .A(images_bus[440]), .ZN(n9484) );
  oai21d1 U5495 ( .B1(n4301), .B2(n3111), .A(n3090), .ZN(n9482) );
  oai211d1 U5497 ( .C1(n9491), .C2(n9492), .A(n9493), .B(n9494), .ZN(n9481) );
  aoi22d1 U5498 ( .A1(n9491), .A2(n6428), .B1(n8736), .B2(n3105), .ZN(n9494)
         );
  aon211d1 U5499 ( .C1(n3014), .C2(n9496), .B(n6428), .A(n7973), .ZN(n9493) );
  aon211d1 U5500 ( .C1(n9497), .C2(n6083), .B(n9498), .A(n2927), .ZN(n9492) );
  aoi31d1 U5502 ( .B1(n9502), .B2(n9503), .B3(n3007), .A(n9501), .ZN(n9499) );
  oai322d1 U5503 ( .C1(n9504), .C2(images_bus[453]), .C3(n3006), .A1(n9506), 
        .A2(n2941), .B1(n6598), .B2(n4792), .ZN(n9503) );
  aoi31d1 U5504 ( .B1(n3004), .B2(n9508), .B3(n4798), .A(n9509), .ZN(n9506) );
  oan211d1 U5505 ( .C1(n8047), .C2(n9510), .B(n9511), .A(n9512), .ZN(n9509) );
  aor31d1 U5506 ( .B1(n2956), .B2(n9514), .B3(n4814), .A(n9515), .Z(n9508) );
  oai222d1 U5508 ( .A1(n9516), .A2(n7336), .B1(n9517), .B2(n9518), .C1(
        images_bus[460]), .C2(n3001), .ZN(n9514) );
  oaim21d1 U5509 ( .B1(N14850), .B2(n2994), .A(n6555), .ZN(n9518) );
  aoi311d1 U5510 ( .C1(n8766), .C2(n8767), .C3(n2998), .A(n9521), .B(n8760), 
        .ZN(n9516) );
  oan211d1 U5511 ( .C1(images_bus[463]), .C2(n8769), .B(n9522), .A(n9523), 
        .ZN(n9521) );
  oai321d1 U5514 ( .C1(n9526), .C2(images_bus[469]), .C3(n2973), .B1(n9528), 
        .B2(n9529), .A(n9530), .ZN(n9524) );
  aoi22d1 U5515 ( .A1(n9531), .A2(n7333), .B1(n9528), .B2(n12147), .ZN(n9530)
         );
  oai21d1 U5516 ( .B1(n4299), .B2(n9528), .A(n6512), .ZN(n9531) );
  aon211d1 U5517 ( .C1(n9533), .C2(n5798), .B(n9534), .A(n2974), .ZN(n9529) );
  oan211d1 U5518 ( .C1(n9535), .C2(n9536), .B(n9537), .A(n9538), .ZN(n9534) );
  aoi31d1 U5520 ( .B1(n4850), .B2(n12151), .B3(n2982), .A(n9541), .ZN(n9535)
         );
  aoi211d1 U5521 ( .C1(images_bus[477]), .C2(n9542), .A(n9543), .B(n9544), 
        .ZN(n9541) );
  oan211d1 U5522 ( .C1(n9545), .C2(n9546), .B(n9547), .A(n9542), .ZN(n9544) );
  oan211d1 U5524 ( .C1(images_bus[484]), .C2(n9548), .B(n9549), .A(n2848), 
        .ZN(n9546) );
  aon211d1 U5526 ( .C1(n8802), .C2(n9552), .B(n2857), .A(n9554), .ZN(n9549) );
  oai211d1 U5528 ( .C1(n7341), .C2(n2862), .A(n9557), .B(n9558), .ZN(n9552) );
  aon211d1 U5529 ( .C1(n2877), .C2(n9559), .B(n9560), .A(n8005), .ZN(n9558) );
  oai322d1 U5531 ( .C1(n9562), .C2(images_bus[493]), .C3(n9563), .A1(n9564), 
        .A2(n9565), .B1(images_bus[492]), .B2(n2872), .ZN(n9559) );
  aoi321d1 U5532 ( .C1(n2878), .C2(n9568), .C3(n2884), .B1(n8810), .B2(n8815), 
        .A(n9569), .ZN(n9564) );
  aoi211d1 U5533 ( .C1(n8811), .C2(n8820), .A(n8810), .B(images_bus[495]), 
        .ZN(n9569) );
  oai321d1 U5534 ( .C1(n8016), .C2(n9570), .C3(n2891), .B1(images_bus[500]), 
        .B2(n9571), .A(n9572), .ZN(n9568) );
  aoi22d1 U5536 ( .A1(n2903), .A2(n9573), .B1(n8026), .B2(n9574), .ZN(n9571)
         );
  aoi322d1 U5537 ( .C1(n2896), .C2(n9576), .C3(n9577), .A1(n9578), .A2(n9579), 
        .B1(n9580), .B2(n5797), .ZN(n9570) );
  aor22d1 U5538 ( .A1(n9581), .A2(n2889), .B1(n9577), .B2(n9583), .Z(n9580) );
  oai21d1 U5539 ( .B1(n6423), .B2(n2898), .A(n8826), .ZN(n9576) );
  aon211d1 U5541 ( .C1(n2862), .C2(n9584), .B(n9585), .A(n5968), .ZN(n9557) );
  aoi31d1 U5543 ( .B1(n2864), .B2(n9590), .B3(n9591), .A(n9592), .ZN(n9548) );
  aoi211d1 U5544 ( .C1(n2859), .C2(n2864), .A(n9594), .B(n2912), .ZN(n9592) );
  aoi22d1 U5545 ( .A1(n2847), .A2(n8787), .B1(images_bus[479]), .B2(n2914), 
        .ZN(n9545) );
  aoi31d1 U5546 ( .B1(images_bus[465]), .B2(n9597), .B3(images_bus[464]), .A(
        n9598), .ZN(n8769) );
  oan211d1 U5548 ( .C1(n3094), .C2(n4300), .B(n9599), .A(n6519), .ZN(n9478) );
  oai21d1 U5550 ( .B1(n3079), .B2(n8720), .A(n8712), .ZN(n6568) );
  oai22d1 U5555 ( .A1(images_bus[407]), .A2(n9604), .B1(n4303), .B2(n3232), 
        .ZN(n9442) );
  oai21d1 U5557 ( .B1(n4970), .B2(n9406), .A(n4968), .ZN(n9416) );
  aoi21d1 U5562 ( .B1(images_bus[371]), .B2(n9397), .A(n6525), .ZN(n9399) );
  aoi21d1 U5565 ( .B1(n6594), .B2(n9607), .A(n3138), .ZN(n8841) );
  aoim21d1 U5571 ( .B1(n5249), .B2(n9377), .A(n12138), .ZN(n9381) );
  oai21d1 U5583 ( .B1(n5046), .B2(n9352), .A(images_bus[340]), .ZN(n9356) );
  or02d0 U5585 ( .A1(n9349), .A2(n5927), .Z(n9347) );
  oai21d1 U5593 ( .B1(n5254), .B2(n9328), .A(images_bus[324]), .ZN(n9331) );
  aoim21d1 U5602 ( .B1(n4939), .B2(n9314), .A(n6455), .ZN(n9320) );
  aoi21d1 U5609 ( .B1(images_bus[307]), .B2(n9298), .A(n12146), .ZN(n9302) );
  aoi31d1 U5610 ( .B1(images_bus[303]), .B2(n4439), .B3(n9292), .A(n5535), 
        .ZN(n9298) );
  oai21d1 U5611 ( .B1(n4439), .B2(n7078), .A(n9292), .ZN(n9295) );
  aoi31d1 U5612 ( .B1(images_bus[296]), .B2(n9290), .B3(n5165), .A(n6565), 
        .ZN(n9292) );
  aoi21d1 U5615 ( .B1(images_bus[291]), .B2(n3493), .A(n6613), .ZN(n9283) );
  aoi21d1 U5622 ( .B1(n4946), .B2(n9264), .A(n12149), .ZN(n9267) );
  aoim21d1 U5623 ( .B1(n5834), .B2(n9256), .A(n6612), .ZN(n9264) );
  oai311d1 U5625 ( .C1(n5740), .C2(n9618), .C3(n5060), .A(images_bus[276]), 
        .B(n9619), .ZN(n9256) );
  aoi211d1 U5626 ( .C1(n9251), .C2(images_bus[267]), .A(n7406), .B(n6566), 
        .ZN(n9618) );
  oaim311d1 U5631 ( .C1(n4442), .C2(n9238), .C3(images_bus[259]), .A(n9621), 
        .B(n6134), .ZN(n9244) );
  oai21d1 U5637 ( .B1(n5063), .B2(n9216), .A(images_bus[244]), .ZN(n9219) );
  oai211d1 U5639 ( .C1(n8078), .C2(n3717), .A(images_bus[240]), .B(n5544), 
        .ZN(n9216) );
  aoi21d1 U5641 ( .B1(images_bus[235]), .B2(n9211), .A(n6567), .ZN(n9214) );
  aoi21d1 U5650 ( .B1(images_bus[227]), .B2(n9191), .A(n12137), .ZN(n9193) );
  ora311d1 U5651 ( .C1(n9181), .C2(n6115), .C3(n7711), .A(images_bus[224]), 
        .B(n5748), .Z(n9191) );
  aor31d1 U5652 ( .B1(n8421), .B2(n9178), .B3(images_bus[216]), .A(n6475), .Z(
        n9181) );
  aoi21d1 U5655 ( .B1(images_bus[211]), .B2(n9173), .A(n6540), .ZN(n9176) );
  aoi21d1 U5667 ( .B1(n9151), .B2(n7422), .A(n6628), .ZN(n9154) );
  oai21d1 U5669 ( .B1(n12168), .B2(n9149), .A(images_bus[188]), .ZN(n9145) );
  aoi31d1 U5679 ( .B1(images_bus[171]), .B2(n9128), .B3(n8866), .A(n6572), 
        .ZN(n9129) );
  oai211d1 U5686 ( .C1(n3982), .C2(n9119), .A(images_bus[163]), .B(n5780), 
        .ZN(n9634) );
  oai31d1 U5687 ( .B1(n4959), .B2(n9113), .B3(n7434), .A(images_bus[156]), 
        .ZN(n9119) );
  aoi21d1 U5690 ( .B1(images_bus[147]), .B2(n9108), .A(n12144), .ZN(n9115) );
  aoi21d1 U5691 ( .B1(n4471), .B2(n9102), .A(n9636), .ZN(n9108) );
  oai21d1 U5699 ( .B1(n5281), .B2(n9086), .A(n4742), .ZN(n9092) );
  oai21d1 U5700 ( .B1(images_bus[133]), .B2(n9638), .A(images_bus[132]), .ZN(
        n5056) );
  aor21d1 U5701 ( .B1(n3991), .B2(n9078), .A(n5053), .Z(n9086) );
  aoi31d1 U5705 ( .B1(images_bus[123]), .B2(n9077), .B3(n6651), .A(n6488), 
        .ZN(n9078) );
  aoi21d1 U5707 ( .B1(images_bus[115]), .B2(n9063), .A(n12143), .ZN(n9069) );
  aoi211d1 U5708 ( .C1(n7440), .C2(n4137), .A(n7097), .B(n5926), .ZN(n9063) );
  aoim21d1 U5713 ( .B1(n5284), .B2(n9035), .A(n6639), .ZN(n9042) );
  oai211d1 U5714 ( .C1(n4139), .C2(n9031), .A(images_bus[96]), .B(n5890), .ZN(
        n9035) );
  aoi21d1 U5718 ( .B1(images_bus[83]), .B2(n9020), .A(n6548), .ZN(n9023) );
  aoi311d1 U5719 ( .C1(n4142), .C2(n4510), .C3(images_bus[79]), .A(n7104), .B(
        n6662), .ZN(n9020) );
  oai21d1 U5721 ( .B1(n5204), .B2(n9013), .A(images_bus[76]), .ZN(n9015) );
  nd13d1 U5722 ( .A1(n9010), .A2(images_bus[72]), .A3(n5693), .ZN(n9013) );
  or02d0 U5724 ( .A1(n8996), .A2(n5815), .Z(n9007) );
  oai21d1 U5725 ( .B1(n5298), .B2(n8993), .A(images_bus[68]), .ZN(n8996) );
  aoi31d1 U5728 ( .B1(n5465), .B2(n4283), .B3(images_bus[59]), .A(n6502), .ZN(
        n8984) );
  oai21d1 U5734 ( .B1(n5110), .B2(n8959), .A(images_bus[52]), .ZN(n8970) );
  oaim21d1 U5735 ( .B1(n6719), .B2(n4285), .A(n7456), .ZN(n8959) );
  oai21d1 U5737 ( .B1(n5205), .B2(n8948), .A(images_bus[44]), .ZN(n8951) );
  or04d0 U5738 ( .A1(n5704), .A2(n7183), .A3(n6884), .A4(n8946), .Z(n8948) );
  aoi21d1 U5742 ( .B1(n9643), .B2(n6688), .A(n6646), .ZN(n8936) );
  aoi31d1 U5743 ( .B1(images_bus[31]), .B2(n8126), .B3(n8933), .A(n5312), .ZN(
        n9643) );
  aoi31d1 U5744 ( .B1(images_bus[24]), .B2(n8926), .B3(n8127), .A(n6507), .ZN(
        n8933) );
  aoi31d1 U5746 ( .B1(images_bus[19]), .B2(n4530), .B3(n5595), .A(n6552), .ZN(
        n8921) );
  oai21d1 U5751 ( .B1(n4866), .B2(n8141), .A(images_bus[12]), .ZN(n8907) );
  oai21d1 U5757 ( .B1(n9645), .B2(n2773), .A(n9647), .ZN(N26359) );
  aor211d1 U5758 ( .C1(n2810), .C2(n9649), .A(n8130), .B(n7461), .Z(n9647) );
  oan211d1 U5762 ( .C1(n9654), .C2(n4771), .B(n9656), .A(n9657), .ZN(n9653) );
  aoi321d1 U5763 ( .C1(n7466), .C2(n9658), .C3(n9659), .B1(n4793), .B2(n5220), 
        .A(n9660), .ZN(n9654) );
  oai221d1 U5765 ( .B1(n9662), .B2(n7462), .C1(n9663), .C2(n9664), .A(n9665), 
        .ZN(n9658) );
  aoi22d1 U5766 ( .A1(n9666), .A2(n7468), .B1(n9667), .B2(n4587), .ZN(n9662)
         );
  oan211d1 U5767 ( .C1(n4619), .C2(n9670), .B(images_bus[18]), .A(n9671), .ZN(
        n9667) );
  oan211d1 U5768 ( .C1(n4619), .C2(n6552), .B(n9672), .A(n8888), .ZN(n9666) );
  aon211d1 U5769 ( .C1(n4365), .C2(n4352), .B(n9675), .A(n4576), .ZN(n9672) );
  aoi31d1 U5770 ( .B1(n9677), .B2(images_bus[23]), .B3(n9678), .A(n9679), .ZN(
        n9675) );
  oan211d1 U5771 ( .C1(n9680), .C2(n9681), .B(n4368), .A(n4366), .ZN(n9678) );
  aoi311d1 U5777 ( .C1(n4347), .C2(images_bus[27]), .C3(n9686), .A(n9687), .B(
        n9688), .ZN(n9680) );
  aoi21d1 U5778 ( .B1(n4376), .B2(n9689), .A(n9690), .ZN(n9686) );
  oai22d1 U5779 ( .A1(images_bus[30]), .A2(n9691), .B1(n9692), .B2(n6671), 
        .ZN(n9689) );
  aoi211d1 U5780 ( .C1(n4232), .C2(n9694), .A(n9695), .B(n7498), .ZN(n9692) );
  oai211d1 U5782 ( .C1(n9699), .C2(n4238), .A(n9700), .B(n9701), .ZN(n9694) );
  aoi211d1 U5783 ( .C1(n7500), .C2(n9702), .A(n9703), .B(n4246), .ZN(n9699) );
  oai211d1 U5785 ( .C1(n9705), .C2(n5800), .A(n9706), .B(n9707), .ZN(n9702) );
  aon211d1 U5786 ( .C1(n4273), .C2(n9708), .B(n6884), .A(n4272), .ZN(n9707) );
  aoi311d1 U5787 ( .C1(n6720), .C2(n9710), .C3(n5789), .A(n9711), .B(n9712), 
        .ZN(n9705) );
  oan211d1 U5788 ( .C1(n9713), .C2(n8957), .B(images_bus[46]), .A(n6713), .ZN(
        n9711) );
  oai222d1 U5790 ( .A1(n9715), .A2(n4252), .B1(n9717), .B2(n9718), .C1(n9719), 
        .C2(n4255), .ZN(n9710) );
  aoi21d1 U5791 ( .B1(n8967), .B2(n9720), .A(n9721), .ZN(n9717) );
  aoi31d1 U5792 ( .B1(images_bus[55]), .B2(n9722), .B3(n4225), .A(n8974), .ZN(
        n9721) );
  oai311d1 U5795 ( .C1(n8116), .C2(n9728), .C3(n8992), .A(n9729), .B(n9730), 
        .ZN(n9727) );
  aoi21d1 U5796 ( .B1(n9731), .B2(n9732), .A(n6701), .ZN(n9730) );
  aoi31d1 U5797 ( .B1(n9733), .B2(n8988), .B3(n9734), .A(n9735), .ZN(n9728) );
  oan211d1 U5798 ( .C1(n9736), .C2(n9737), .B(n9738), .A(n4222), .ZN(n9734) );
  aoi31d1 U5799 ( .B1(n5033), .B2(n4186), .B3(n9740), .A(n9741), .ZN(n9736) );
  aoi21d1 U5800 ( .B1(n9742), .B2(n9743), .A(n5793), .ZN(n9741) );
  aoi22d1 U5801 ( .A1(n6744), .A2(n9744), .B1(n4189), .B2(n9745), .ZN(n9742)
         );
  oan211d1 U5803 ( .C1(n9747), .C2(n5020), .B(n9748), .A(n5793), .ZN(n9740) );
  aoi311d1 U5804 ( .C1(n4180), .C2(n9749), .C3(n4151), .A(n9751), .B(n9752), 
        .ZN(n9747) );
  oan211d1 U5805 ( .C1(n9753), .C2(n8112), .B(images_bus[74]), .A(n9012), .ZN(
        n9751) );
  oai22d1 U5806 ( .A1(n9753), .A2(n6586), .B1(n9754), .B2(n4155), .ZN(n9749)
         );
  aoi221d1 U5807 ( .B1(n7548), .B2(n9755), .C1(n4178), .C2(n4223), .A(n9757), 
        .ZN(n9754) );
  oai322d1 U5809 ( .C1(n9759), .C2(n4161), .C3(n9761), .A1(n9762), .A2(n5848), 
        .B1(n9758), .B2(n7104), .ZN(n9755) );
  aoi321d1 U5810 ( .C1(n7557), .C2(n9763), .C3(n4173), .B1(n4175), .B2(n5106), 
        .A(n9764), .ZN(n9762) );
  oai211d1 U5811 ( .C1(n9765), .C2(n5858), .A(n4172), .B(n4176), .ZN(n9759) );
  aoi211d1 U5812 ( .C1(n9767), .C2(n9768), .A(n5866), .B(n9769), .ZN(n9765) );
  aoi31d1 U5814 ( .B1(n9767), .B2(images_bus[91]), .B3(n9772), .A(n7447), .ZN(
        n9771) );
  aoi311d1 U5815 ( .C1(n4117), .C2(n4170), .C3(n9773), .A(n9774), .B(n9775), 
        .ZN(n9772) );
  oan211d1 U5817 ( .C1(n9778), .C2(n5884), .B(n9779), .A(n9777), .ZN(n9773) );
  aoi221d1 U5819 ( .B1(n4112), .B2(n9781), .C1(n4116), .C2(n9782), .A(n9783), 
        .ZN(n9778) );
  oai311d1 U5820 ( .C1(n7573), .C2(n9784), .C3(n7176), .A(n9785), .B(n5885), 
        .ZN(n9783) );
  aoi221d1 U5822 ( .B1(images_bus[104]), .B2(n9786), .C1(n4072), .C2(n9788), 
        .A(n9789), .ZN(n9784) );
  aoi21d1 U5823 ( .B1(n9790), .B2(n6799), .A(n9791), .ZN(n9789) );
  oai211d1 U5824 ( .C1(n9792), .C2(n5917), .A(n9062), .B(n9793), .ZN(n9788) );
  oai21d1 U5825 ( .B1(n5203), .B2(n4060), .A(images_bus[108]), .ZN(n9793) );
  aoi31d1 U5828 ( .B1(n4081), .B2(n4108), .B3(n9796), .A(n9797), .ZN(n9792) );
  aoi31d1 U5829 ( .B1(n9798), .B2(n9799), .B3(n4058), .A(n7583), .ZN(n9796) );
  aon211d1 U5831 ( .C1(n4099), .C2(n9803), .B(n4059), .A(n5036), .ZN(n9798) );
  oai211d1 U5832 ( .C1(n9805), .C2(n4089), .A(n7439), .B(n9807), .ZN(n9803) );
  aoi22d1 U5834 ( .A1(n4092), .A2(n9809), .B1(n4091), .B2(n4965), .ZN(n9805)
         );
  oai31d1 U5836 ( .B1(n5040), .B2(n9810), .B3(n9811), .A(n9812), .ZN(n9809) );
  aoi211d1 U5837 ( .C1(n8307), .C2(n9813), .A(n9814), .B(n9815), .ZN(n9810) );
  oai22d1 U5838 ( .A1(images_bus[126]), .A2(n5951), .B1(n9816), .B2(n5041), 
        .ZN(n9814) );
  oai211d1 U5839 ( .C1(n9817), .C2(n5050), .A(n9818), .B(n9819), .ZN(n9813) );
  aoi22d1 U5840 ( .A1(n5771), .A2(n3985), .B1(n4006), .B2(n6946), .ZN(n9819)
         );
  oai321d1 U5842 ( .C1(n8320), .C2(n9823), .C3(n8322), .B1(n9824), .B2(n4016), 
        .A(n9825), .ZN(n9822) );
  aoi21d1 U5843 ( .B1(n9098), .B2(n9826), .A(n9827), .ZN(n9825) );
  aoi31d1 U5846 ( .B1(n7620), .B2(n4024), .B3(n9829), .A(n5194), .ZN(n9824) );
  aoi22d1 U5847 ( .A1(n9830), .A2(n9831), .B1(n9832), .B2(n5076), .ZN(n9829)
         );
  aon211d1 U5848 ( .C1(n4051), .C2(n9833), .B(n9834), .A(n4027), .ZN(n9831) );
  oai22d1 U5849 ( .A1(n9835), .A2(n9836), .B1(n9837), .B2(n5095), .ZN(n9833)
         );
  oai211d1 U5851 ( .C1(n7644), .C2(n9841), .A(n9842), .B(n9843), .ZN(n9838) );
  aoi21d1 U5852 ( .B1(n4033), .B2(n9844), .A(n9845), .ZN(n9843) );
  oai22d1 U5853 ( .A1(images_bus[154]), .A2(n8337), .B1(n9846), .B2(n9847), 
        .ZN(n9844) );
  aon211d1 U5854 ( .C1(n9848), .C2(n6185), .B(n9849), .A(n4043), .ZN(n9841) );
  aon211d1 U5855 ( .C1(n9850), .C2(n9851), .B(n5984), .A(n3902), .ZN(n9849) );
  oai211d1 U5858 ( .C1(n9855), .C2(n9856), .A(n9857), .B(n3911), .ZN(n9851) );
  oai22d1 U5859 ( .A1(n9858), .A2(n6880), .B1(n9859), .B2(n9860), .ZN(n9856)
         );
  aoi211d1 U5861 ( .C1(n3922), .C2(n9862), .A(n9863), .B(n9864), .ZN(n9858) );
  aoi211d1 U5864 ( .C1(n3929), .C2(n9868), .A(n9869), .B(n6866), .ZN(n9865) );
  aon211d1 U5865 ( .C1(n9870), .C2(n9871), .B(n9872), .A(n9873), .ZN(n9869) );
  aon211d1 U5866 ( .C1(n9632), .C2(n9874), .B(n9875), .A(n9876), .ZN(n9871) );
  oai211d1 U5867 ( .C1(n9877), .C2(n3940), .A(n9879), .B(n9880), .ZN(n9874) );
  aoi311d1 U5871 ( .C1(n3962), .C2(n9881), .C3(n3950), .A(n9882), .B(n9883), 
        .ZN(n9877) );
  oai22d1 U5872 ( .A1(images_bus[182]), .A2(n7428), .B1(n9884), .B2(n3946), 
        .ZN(n9882) );
  oai222d1 U5875 ( .A1(n9885), .A2(n6927), .B1(n9884), .B2(n9886), .C1(n9887), 
        .C2(n3959), .ZN(n9881) );
  aoi21d1 U5876 ( .B1(n3957), .B2(n9888), .A(n9889), .ZN(n9885) );
  oai222d1 U5877 ( .A1(n9887), .A2(n6481), .B1(n9890), .B2(n5187), .C1(n9891), 
        .C2(n9892), .ZN(n9888) );
  aoi21d1 U5878 ( .B1(n6013), .B2(n9893), .A(n9894), .ZN(n9890) );
  oai22d1 U5879 ( .A1(n9895), .A2(n9896), .B1(n9897), .B2(n4390), .ZN(n9893)
         );
  aoi311d1 U5880 ( .C1(n3834), .C2(n3880), .C3(n9898), .A(n3812), .B(n5276), 
        .ZN(n9897) );
  aoi31d1 U5881 ( .B1(n9900), .B2(n9901), .B3(n9902), .A(n9903), .ZN(n9898) );
  aoi21d1 U5882 ( .B1(n3836), .B2(n9904), .A(n6390), .ZN(n9902) );
  aon211d1 U5883 ( .C1(n3844), .C2(n12128), .B(n9906), .A(n6031), .ZN(n9900)
         );
  oan211d1 U5884 ( .C1(n9907), .C2(n6943), .B(n9908), .A(n5209), .ZN(n9906) );
  oai321d1 U5887 ( .C1(n9910), .C2(n9911), .C3(n5230), .B1(n3811), .B2(n5227), 
        .A(n9913), .ZN(n9909) );
  or02d0 U5889 ( .A1(n5227), .A2(n4388), .Z(n5230) );
  aor31d1 U5890 ( .B1(n5236), .B2(n9915), .B3(n9916), .A(n5548), .Z(n9910) );
  aoi22d1 U5891 ( .A1(n9917), .A2(n3851), .B1(n3875), .B2(n9918), .ZN(n9916)
         );
  aoi31d1 U5893 ( .B1(n9920), .B2(n9921), .B3(n9922), .A(n5244), .ZN(n9917) );
  aoi22d1 U5894 ( .A1(n3868), .A2(n9923), .B1(n5240), .B2(n6250), .ZN(n9922)
         );
  oai321d1 U5896 ( .C1(n9185), .C2(n9927), .C3(n6059), .B1(n9928), .B2(n9929), 
        .A(n9930), .ZN(n9926) );
  aoim211d1 U5897 ( .C1(n5270), .C2(n3736), .A(n9931), .B(n9932), .ZN(n9927)
         );
  oan211d1 U5898 ( .C1(n9933), .C2(n3730), .B(n9934), .A(n9935), .ZN(n9932) );
  aoi211d1 U5899 ( .C1(n3742), .C2(n5268), .A(n9936), .B(n9937), .ZN(n9933) );
  oan211d1 U5900 ( .C1(n9938), .C2(n9939), .B(images_bus[230]), .A(n9940), 
        .ZN(n9937) );
  aoi211d1 U5901 ( .C1(n3757), .C2(n9941), .A(n9942), .B(n6389), .ZN(n9938) );
  aon211d1 U5902 ( .C1(n9943), .C2(n9944), .B(n3755), .A(n9946), .ZN(n9942) );
  oan211d1 U5905 ( .C1(n9947), .C2(n9948), .B(n7724), .A(n9949), .ZN(n9943) );
  oai22d1 U5908 ( .A1(n9950), .A2(n8445), .B1(n9951), .B2(n8442), .ZN(n9948)
         );
  oai211d1 U5909 ( .C1(n9952), .C2(n9953), .A(n3770), .B(n3801), .ZN(n8442) );
  oai22d1 U5911 ( .A1(n9954), .A2(n9955), .B1(n9956), .B2(n8449), .ZN(n9947)
         );
  aoi22d1 U5914 ( .A1(n3795), .A2(n9959), .B1(images_bus[244]), .B2(n9960), 
        .ZN(n9956) );
  oai221d1 U5915 ( .B1(n9961), .B2(n3781), .C1(n3586), .C2(n9227), .A(n9963), 
        .ZN(n9959) );
  aoi221d1 U5918 ( .B1(n6111), .B2(n4948), .C1(images_bus[248]), .C2(n9964), 
        .A(n9965), .ZN(n9961) );
  oan211d1 U5919 ( .C1(n9966), .C2(n4410), .B(n9967), .A(n7011), .ZN(n9965) );
  aoi31d1 U5923 ( .B1(images_bus[254]), .B2(n9971), .B3(n9972), .A(n5347), 
        .ZN(n9969) );
  aoi31d1 U5924 ( .B1(n3570), .B2(n5266), .B3(n7027), .A(n9974), .ZN(n9972) );
  aoi321d1 U5927 ( .C1(n9977), .C2(n9978), .C3(n3531), .B1(n8471), .B2(n6024), 
        .A(n3505), .ZN(n9975) );
  oai22d1 U5930 ( .A1(images_bus[263]), .A2(n9982), .B1(n9983), .B2(n7031), 
        .ZN(n9978) );
  aoi221d1 U5931 ( .B1(n5745), .B2(n9984), .C1(n3566), .C2(n9986), .A(n9987), 
        .ZN(n9983) );
  oai322d1 U5932 ( .C1(n7037), .C2(n9988), .C3(n9989), .A1(n9990), .A2(n6616), 
        .B1(images_bus[270]), .B2(n7760), .ZN(n9984) );
  aoi22d1 U5933 ( .A1(n7040), .A2(n9991), .B1(images_bus[272]), .B2(n3507), 
        .ZN(n9988) );
  aon211d1 U5934 ( .C1(n9993), .C2(n9994), .B(n7041), .A(n9995), .ZN(n9991) );
  aon211d1 U5935 ( .C1(n3540), .C2(n5060), .B(n3506), .A(n9998), .ZN(n9995) );
  oan211d1 U5938 ( .C1(n10000), .C2(n10001), .B(n7035), .A(n10002), .ZN(n9994)
         );
  aoi21d1 U5939 ( .B1(n9999), .B2(images_bus[275]), .A(n6533), .ZN(n10002) );
  aoi31d1 U5942 ( .B1(n10004), .B2(n4946), .B3(n10005), .A(n7044), .ZN(n10000)
         );
  aon211d1 U5943 ( .C1(n7046), .C2(n10006), .B(n6173), .A(n3476), .ZN(n10005)
         );
  oai211d1 U5945 ( .C1(n10007), .C2(n9273), .A(images_bus[286]), .B(n10008), 
        .ZN(n10006) );
  aoi21d1 U5946 ( .B1(n3423), .B2(n10009), .A(n3484), .ZN(n10008) );
  aon211d1 U5947 ( .C1(n10011), .C2(n10012), .B(n10013), .A(n10014), .ZN(
        n10009) );
  aoi21d1 U5948 ( .B1(n3428), .B2(n10015), .A(n10016), .ZN(n10011) );
  oai322d1 U5949 ( .C1(n4495), .C2(n10017), .C3(n5396), .A1(n10018), .A2(n9289), .B1(n6383), .B2(n5392), .ZN(n10015) );
  oai211d1 U5950 ( .C1(n10019), .C2(n10020), .A(n3469), .B(n3471), .ZN(n9289)
         );
  aoi221d1 U5952 ( .B1(n3466), .B2(n6842), .C1(n3464), .C2(n10021), .A(n10022), 
        .ZN(n10017) );
  oai31d1 U5953 ( .B1(n10023), .B2(n10024), .B3(n5402), .A(n10025), .ZN(n10021) );
  aoi221d1 U5954 ( .B1(images_bus[300]), .B2(n3483), .C1(n3432), .C2(n10027), 
        .A(n10028), .ZN(n10024) );
  oan211d1 U5955 ( .C1(n10029), .C2(n8526), .B(n10030), .A(n7078), .ZN(n10028)
         );
  oai22d1 U5956 ( .A1(n10031), .A2(n5403), .B1(n10032), .B2(n9303), .ZN(n10027) );
  aoi311d1 U5957 ( .C1(n3451), .C2(n3458), .C3(n10033), .A(n5049), .B(n10034), 
        .ZN(n10032) );
  oan211d1 U5959 ( .C1(n10036), .C2(n3441), .B(n10038), .A(n5049), .ZN(n10033)
         );
  aoi211d1 U5962 ( .C1(n3443), .C2(n10040), .A(n10041), .B(n10042), .ZN(n10036) );
  aoi21d1 U5963 ( .B1(n3482), .B2(n10044), .A(n10045), .ZN(n10042) );
  oai211d1 U5964 ( .C1(n10046), .C2(n10047), .A(n3420), .B(n6194), .ZN(n10044)
         );
  oan211d1 U5966 ( .C1(n10049), .C2(n10050), .B(n10051), .A(n6198), .ZN(n10046) );
  aon211d1 U5967 ( .C1(n3364), .C2(n3333), .B(n10053), .A(n10054), .ZN(n10050)
         );
  aoi311d1 U5968 ( .C1(n10055), .C2(n6204), .C3(n10056), .A(n10057), .B(n6197), 
        .ZN(n10053) );
  aon211d1 U5969 ( .C1(n10058), .C2(n3416), .B(n10059), .A(n3367), .ZN(n10055)
         );
  aoi31d1 U5970 ( .B1(n10060), .B2(n10061), .B3(n10062), .A(n4545), .ZN(n10059) );
  aoi22d1 U5971 ( .A1(n4548), .A2(n10063), .B1(n3411), .B2(n10064), .ZN(n10062) );
  oai322d1 U5973 ( .C1(n5445), .C2(n10066), .C3(n10067), .A1(n3332), .A2(n7136), .B1(n10069), .B2(n3407), .ZN(n10065) );
  aoi311d1 U5976 ( .C1(n3377), .C2(n10072), .C3(n3374), .A(n10074), .B(n10075), 
        .ZN(n10066) );
  aoi21d1 U5977 ( .B1(n10076), .B2(images_bus[335]), .A(n10077), .ZN(n10075)
         );
  oaim22d1 U5978 ( .A1(n10076), .A2(n7123), .B1(n10063), .B2(images_bus[332]), 
        .ZN(n10074) );
  aoi31d1 U5979 ( .B1(images_bus[333]), .B2(n10063), .B3(images_bus[332]), .A(
        n6297), .ZN(n10076) );
  aoi31d1 U5981 ( .B1(images_bus[329]), .B2(n10064), .B3(images_bus[328]), .A(
        n6840), .ZN(n10069) );
  oai211d1 U5984 ( .C1(images_bus[339]), .C2(n6252), .A(n10078), .B(
        images_bus[338]), .ZN(n10072) );
  aon211d1 U5985 ( .C1(n3398), .C2(n12157), .B(n10079), .A(n7135), .ZN(n10078)
         );
  oan211d1 U5986 ( .C1(n7139), .C2(n10080), .B(images_bus[343]), .A(n10081), 
        .ZN(n10079) );
  aon211d1 U5987 ( .C1(n10082), .C2(n8581), .B(n10083), .A(n3395), .ZN(n10080)
         );
  aoi22d1 U5988 ( .A1(images_bus[347]), .A2(images_bus[346]), .B1(
        images_bus[346]), .B2(n8570), .ZN(n10083) );
  oan211d1 U5989 ( .C1(n10085), .C2(n10086), .B(images_bus[350]), .A(n3391), 
        .ZN(n10082) );
  oan211d1 U5990 ( .C1(n10087), .C2(n10088), .B(n7850), .A(n6097), .ZN(n10085)
         );
  oai22d1 U5993 ( .A1(images_bus[355]), .A2(n10090), .B1(n10091), .B2(n5478), 
        .ZN(n10088) );
  aoi22d1 U5995 ( .A1(n3318), .A2(n5988), .B1(n6299), .B2(n10093), .ZN(n10091)
         );
  oai221d1 U5996 ( .B1(images_bus[363]), .B2(n7381), .C1(n10094), .C2(n4602), 
        .A(images_bus[362]), .ZN(n10093) );
  aoi31d1 U5997 ( .B1(n3313), .B2(n10096), .B3(n6316), .A(n5146), .ZN(n10094)
         );
  oai211d1 U5998 ( .C1(images_bus[367]), .C2(n10097), .A(n10098), .B(
        images_bus[366]), .ZN(n10096) );
  aon211d1 U5999 ( .C1(n10099), .C2(n10100), .B(n12132), .A(n3287), .ZN(n10098) );
  aon211d1 U6003 ( .C1(images_bus[371]), .C2(n10103), .B(n4623), .A(n6737), 
        .ZN(n10100) );
  oai211d1 U6004 ( .C1(n6229), .C2(n10104), .A(n7189), .B(n3308), .ZN(n10103)
         );
  oai21d1 U6007 ( .B1(images_bus[375]), .B2(n5500), .A(n10107), .ZN(n10104) );
  oan211d1 U6009 ( .C1(n6664), .C2(n3298), .B(n10111), .A(n5512), .ZN(n10108)
         );
  aon211d1 U6010 ( .C1(n10112), .C2(n6353), .B(n10113), .A(n3298), .ZN(n10111)
         );
  aoi221d1 U6012 ( .B1(n9607), .B2(n6162), .C1(n10115), .C2(n3162), .A(n10117), 
        .ZN(n10114) );
  oan211d1 U6013 ( .C1(n10118), .C2(n3250), .B(n10119), .A(n10120), .ZN(n10117) );
  oai211d1 U6014 ( .C1(n10121), .C2(n10122), .A(n3250), .B(n3248), .ZN(n10119)
         );
  oai21d1 U6015 ( .B1(n10123), .B2(n10124), .A(n10125), .ZN(n10122) );
  aon211d1 U6016 ( .C1(n10126), .C2(n10127), .B(n10128), .A(n3171), .ZN(n10125) );
  oan211d1 U6018 ( .C1(n3187), .C2(n10131), .B(n10132), .A(n7225), .ZN(n10128)
         );
  aon211d1 U6019 ( .C1(n7230), .C2(n10133), .B(n10134), .A(n3187), .ZN(n10132)
         );
  oan211d1 U6020 ( .C1(n7889), .C2(n10135), .B(n3184), .A(n10137), .ZN(n10134)
         );
  oai322d1 U6022 ( .C1(n7236), .C2(images_bus[399]), .C3(n3192), .A1(n7893), 
        .A2(n10140), .B1(n10141), .B2(n10142), .ZN(n10133) );
  aon211d1 U6024 ( .C1(n3240), .C2(n10143), .B(n10144), .A(n3205), .ZN(n10140)
         );
  aoi21d1 U6025 ( .B1(n3240), .B2(n8837), .A(n3139), .ZN(n10144) );
  oai322d1 U6027 ( .C1(n10147), .C2(n9438), .C3(n8649), .A1(n10148), .A2(
        n10149), .B1(images_bus[403]), .B2(n8837), .ZN(n10143) );
  aoi31d1 U6028 ( .B1(n3238), .B2(n8651), .B3(n3207), .A(n8644), .ZN(n10148)
         );
  aon211d1 U6031 ( .C1(n3217), .C2(n10151), .B(n10152), .A(n3211), .ZN(n10147)
         );
  aon211d1 U6032 ( .C1(images_bus[406]), .C2(n10149), .B(n3232), .A(n10153), 
        .ZN(n10152) );
  aon211d1 U6033 ( .C1(n3219), .C2(n10155), .B(n10156), .A(n9447), .ZN(n10153)
         );
  oai31d1 U6034 ( .B1(n8658), .B2(n3222), .B3(n10157), .A(n10158), .ZN(n10156)
         );
  oai211d1 U6036 ( .C1(n10160), .C2(n10161), .A(n10162), .B(n10163), .ZN(
        n10159) );
  aoi31d1 U6037 ( .B1(n10164), .B2(n6577), .B3(n3036), .A(n10166), .ZN(n10163)
         );
  oai21d1 U6041 ( .B1(n10169), .B2(n6160), .A(n8679), .ZN(n10162) );
  aoi31d1 U6042 ( .B1(n6578), .B2(n3133), .B3(images_bus[416]), .A(n10171), 
        .ZN(n10160) );
  oan211d1 U6043 ( .C1(n10172), .C2(n10173), .B(n10174), .A(n3042), .ZN(n10171) );
  aon211d1 U6044 ( .C1(n10176), .C2(n8683), .B(n10177), .A(n10172), .ZN(n10174) );
  aoi211d1 U6045 ( .C1(n8683), .C2(n3127), .A(n10178), .B(n10173), .ZN(n10177)
         );
  oan211d1 U6046 ( .C1(images_bus[421]), .C2(n6448), .B(n6599), .A(n8688), 
        .ZN(n10178) );
  oan211d1 U6047 ( .C1(n3054), .C2(n10179), .B(n10180), .A(n4729), .ZN(n10176)
         );
  aon211d1 U6048 ( .C1(n10181), .C2(n10182), .B(n10183), .A(n3054), .ZN(n10180) );
  aoi21d1 U6049 ( .B1(n9464), .B2(n9469), .A(n10184), .ZN(n10183) );
  oai22d1 U6051 ( .A1(n3123), .A2(n10185), .B1(n10186), .B2(n6460), .ZN(n10182) );
  aoi321d1 U6052 ( .C1(n10187), .C2(n10188), .C3(n10189), .B1(n3068), .B2(
        n10191), .A(n10192), .ZN(n10186) );
  oaim22d1 U6053 ( .A1(n3075), .A2(n10193), .B1(n10194), .B2(n7952), .ZN(
        n10192) );
  oai222d1 U6054 ( .A1(n10195), .A2(n10196), .B1(n10197), .B2(n10198), .C1(
        n6474), .C2(n10199), .ZN(n10191) );
  oaim22d1 U6055 ( .A1(n10200), .A2(n6478), .B1(n6478), .B2(n10201), .ZN(
        n10199) );
  aoi31d1 U6056 ( .B1(n10201), .B2(n6487), .B3(images_bus[438]), .A(n10202), 
        .ZN(n10200) );
  aoi311d1 U6057 ( .C1(n10203), .C2(n10204), .C3(n3110), .A(n6487), .B(n10205), 
        .ZN(n10202) );
  oan211d1 U6058 ( .C1(n10203), .C2(n6990), .B(n3110), .A(n3134), .ZN(n10205)
         );
  oai21d1 U6059 ( .B1(n10207), .B2(n8725), .A(n10208), .ZN(n10204) );
  oai211d1 U6060 ( .C1(n6559), .C2(n7611), .A(n10210), .B(images_bus[440]), 
        .ZN(n10208) );
  aoi322d1 U6063 ( .C1(n10211), .C2(n8726), .C3(n3106), .A1(n10212), .A2(n6557), .B1(n10213), .B2(n3103), .ZN(n10207) );
  oan211d1 U6064 ( .C1(n6428), .C2(n10214), .B(n10215), .A(n6499), .ZN(n10213)
         );
  oai322d1 U6066 ( .C1(n7973), .C2(n10217), .C3(n2936), .A1(n8744), .A2(n10219), .B1(n2927), .B2(n10220), .ZN(n10216) );
  aon211d1 U6067 ( .C1(n10221), .C2(n8030), .B(n10222), .A(n2926), .ZN(n10219)
         );
  oan211d1 U6068 ( .C1(n10223), .C2(n10224), .B(n10225), .A(n8030), .ZN(n10222) );
  oai22d1 U6070 ( .A1(n2951), .A2(n10228), .B1(n10229), .B2(n10230), .ZN(
        n10226) );
  aoi311d1 U6071 ( .C1(n8047), .C2(n7315), .C3(n2918), .A(n10232), .B(n2949), 
        .ZN(n10229) );
  oai22d1 U6073 ( .A1(n10228), .A2(n2948), .B1(n10234), .B2(n2947), .ZN(n10232) );
  aoi211d1 U6075 ( .C1(n2996), .C2(n10237), .A(n10238), .B(n10239), .ZN(n10234) );
  aoi31d1 U6077 ( .B1(n10243), .B2(n6818), .B3(n7316), .A(n10244), .ZN(n10238)
         );
  aoi211d1 U6078 ( .C1(n10245), .C2(n10240), .A(n7316), .B(n10246), .ZN(n10244) );
  aoim21d1 U6079 ( .B1(n7319), .B2(n10247), .A(n10248), .ZN(n10246) );
  aon211d1 U6080 ( .C1(n10249), .C2(n10250), .B(n8766), .A(n10251), .ZN(n10237) );
  oai21d1 U6081 ( .B1(n10245), .B2(n12156), .A(n8766), .ZN(n10251) );
  oai321d1 U6083 ( .C1(n2916), .C2(n10257), .C3(n10258), .B1(n10259), .B2(
        n10260), .A(n10261), .ZN(n10255) );
  aoi21d1 U6084 ( .B1(n10262), .B2(n10258), .A(n10263), .ZN(n10261) );
  aoi31d1 U6085 ( .B1(n10264), .B2(n10265), .B3(n10266), .A(n4837), .ZN(n10263) );
  aoi22d1 U6086 ( .A1(n7987), .A2(n10267), .B1(n4838), .B2(n10268), .ZN(n10266) );
  aon211d1 U6087 ( .C1(n10269), .C2(n10270), .B(n10271), .A(n10272), .ZN(
        n10267) );
  aon211d1 U6088 ( .C1(n9539), .C2(n9536), .B(n9533), .A(n10273), .ZN(n10272)
         );
  oai211d1 U6089 ( .C1(n10274), .C2(n10275), .A(n2982), .B(n2829), .ZN(n10270)
         );
  oan211d1 U6091 ( .C1(n2847), .C2(n10277), .B(n10278), .A(n2845), .ZN(n10274)
         );
  aon211d1 U6094 ( .C1(n10281), .C2(n10282), .B(n10283), .A(n9551), .ZN(n10278) );
  oan211d1 U6096 ( .C1(n10284), .C2(n10285), .B(n10286), .A(n10282), .ZN(
        n10283) );
  oai21d1 U6097 ( .B1(n10285), .B2(n2858), .A(n10281), .ZN(n10286) );
  aoi322d1 U6098 ( .C1(n10288), .C2(n10289), .C3(n8802), .A1(n2858), .A2(n5221), .B1(n2820), .B2(n2863), .ZN(n10284) );
  aon211d1 U6100 ( .C1(images_bus[486]), .C2(n10292), .B(n2862), .A(n10293), 
        .ZN(n10289) );
  aon211d1 U6102 ( .C1(n10297), .C2(n9586), .B(n9584), .A(n10298), .ZN(n10295)
         );
  oan211d1 U6103 ( .C1(n2866), .C2(n10300), .B(n10301), .A(n10297), .ZN(n10294) );
  aoi31d1 U6104 ( .B1(n2871), .B2(n2866), .B3(n10303), .A(n10304), .ZN(n10301)
         );
  oan211d1 U6105 ( .C1(n2821), .C2(n2871), .B(n10306), .A(n10307), .ZN(n10304)
         );
  aon211d1 U6107 ( .C1(n9563), .C2(n2879), .B(n10310), .A(n10311), .ZN(n10309)
         );
  oai322d1 U6109 ( .C1(n8810), .C2(n2822), .C3(n8811), .A1(n10314), .A2(n8813), 
        .B1(images_bus[494]), .B2(n2879), .ZN(n10312) );
  aoi211d1 U6110 ( .C1(n8818), .C2(n10315), .A(n10316), .B(n10317), .ZN(n10314) );
  oan211d1 U6111 ( .C1(n2822), .C2(n8820), .B(n2824), .A(n8821), .ZN(n10317)
         );
  oan211d1 U6113 ( .C1(n4920), .C2(N15458), .B(n2883), .A(n10321), .ZN(n10319)
         );
  oai211d1 U6114 ( .C1(images_bus[497]), .C2(n10322), .A(n4920), .B(
        images_bus[496]), .ZN(n8820) );
  oan211d1 U6115 ( .C1(n4898), .C2(n10323), .B(n10324), .A(n10325), .ZN(n10316) );
  aon211d1 U6116 ( .C1(images_bus[500]), .C2(n10326), .B(n10327), .A(n10328), 
        .ZN(n10324) );
  oai322d1 U6117 ( .C1(n9578), .C2(n10329), .C3(n2823), .A1(n10331), .A2(n4904), .B1(n2889), .B2(n10332), .ZN(n10315) );
  oan211d1 U6118 ( .C1(n9583), .C2(n10333), .B(n10334), .A(n10335), .ZN(n10331) );
  oan211d1 U6119 ( .C1(n2897), .C2(n10337), .B(n10338), .A(n10339), .ZN(n10335) );
  aoi31d1 U6120 ( .B1(n2900), .B2(N15618), .B3(n10341), .A(n10342), .ZN(n10338) );
  aoi211d1 U6121 ( .C1(n10337), .C2(images_bus[507]), .A(n10343), .B(n10344), 
        .ZN(n10342) );
  aoi21d1 U6122 ( .B1(images_bus[509]), .B2(n6423), .A(n2901), .ZN(n10344) );
  aoi31d1 U6124 ( .B1(images_bus[505]), .B2(n10334), .B3(images_bus[504]), .A(
        n6654), .ZN(n10337) );
  aoi31d1 U6131 ( .B1(images_bus[496]), .B2(n10347), .B3(images_bus[497]), .A(
        n6723), .ZN(n10321) );
  aoi21d1 U6134 ( .B1(n8813), .B2(images_bus[496]), .A(n10350), .ZN(n8811) );
  oai211d1 U6137 ( .C1(n5118), .C2(n10351), .A(images_bus[492]), .B(
        images_bus[493]), .ZN(n10310) );
  aoi22d1 U6139 ( .A1(n10352), .A2(n10353), .B1(n2821), .B2(images_bus[491]), 
        .ZN(n10303) );
  oai211d1 U6147 ( .C1(n5221), .C2(n10281), .A(images_bus[484]), .B(
        images_bus[485]), .ZN(n10292) );
  oai21d1 U6148 ( .B1(n10277), .B2(n8830), .A(n6892), .ZN(n10281) );
  aoi31d1 U6150 ( .B1(n10354), .B2(n6425), .B3(images_bus[477]), .A(n12161), 
        .ZN(n10276) );
  oai21d1 U6152 ( .B1(n2913), .B2(n8830), .A(n8832), .ZN(n8029) );
  aon211d1 U6154 ( .C1(n10356), .C2(n6425), .B(n10357), .A(n10354), .ZN(n10269) );
  oaim211d1 U6155 ( .C1(n10273), .C2(n9539), .A(images_bus[474]), .B(
        images_bus[475]), .ZN(n10354) );
  oai21d1 U6157 ( .B1(n4298), .B2(n2916), .A(n6212), .ZN(n10268) );
  oai21d1 U6159 ( .B1(n2831), .B2(n2819), .A(n10359), .ZN(n10356) );
  aon211d1 U6162 ( .C1(images_bus[469]), .C2(n10361), .B(n10362), .A(n10363), 
        .ZN(n10264) );
  aor31d1 U6166 ( .B1(images_bus[464]), .B2(n10364), .B3(images_bus[465]), .A(
        n6731), .Z(n10262) );
  oai21d1 U6168 ( .B1(n10365), .B2(n9598), .A(n10364), .ZN(n10249) );
  aor21d1 U6173 ( .B1(n10366), .B2(images_bus[464]), .A(n10367), .Z(n9598) );
  oaim21d1 U6180 ( .B1(images_bus[455]), .B2(n10228), .A(n8751), .ZN(n10243)
         );
  aoim31d1 U6182 ( .B1(n4635), .B2(n12141), .B3(n10223), .A(n6358), .ZN(n10228) );
  ora31d1 U6183 ( .B1(n2946), .B2(n12141), .B3(n4635), .A(n8746), .Z(n10224)
         );
  oai21d1 U6186 ( .B1(n10217), .B2(n10371), .A(images_bus[450]), .ZN(n10221)
         );
  oai211d1 U6189 ( .C1(n2939), .C2(n10371), .A(n3012), .B(n8050), .ZN(n8740)
         );
  aoim21d1 U6190 ( .B1(n3009), .B2(n10371), .A(n10373), .ZN(n8050) );
  aoi31d1 U6193 ( .B1(images_bus[445]), .B2(n10211), .B3(images_bus[444]), .A(
        n12160), .ZN(n10220) );
  aon211d1 U6194 ( .C1(images_bus[445]), .C2(n8737), .B(n8731), .A(n10211), 
        .ZN(n10214) );
  oai31d1 U6197 ( .B1(n3134), .B2(n12167), .B3(n6990), .A(images_bus[442]), 
        .ZN(n10212) );
  oai211d1 U6200 ( .C1(n5003), .C2(n10375), .A(images_bus[436]), .B(
        images_bus[437]), .ZN(n10201) );
  aoi31d1 U6202 ( .B1(n6563), .B2(n5003), .B3(n3113), .A(n3092), .ZN(n10197)
         );
  oai21d1 U6204 ( .B1(n6563), .B2(n6564), .A(n10375), .ZN(n10378) );
  oai21d1 U6205 ( .B1(n10195), .B2(n8720), .A(images_bus[434]), .ZN(n10375) );
  oai21d1 U6206 ( .B1(n9599), .B2(n6519), .A(n3114), .ZN(n6563) );
  oan211d1 U6209 ( .C1(n3084), .C2(n10382), .B(n3116), .A(n8720), .ZN(n10379)
         );
  aoim31d1 U6218 ( .B1(n5617), .B2(n10184), .B3(n7121), .A(n6826), .ZN(n10185)
         );
  aoim31d1 U6220 ( .B1(n4640), .B2(n12140), .B3(n10173), .A(n6360), .ZN(n10179) );
  oai31d1 U6224 ( .B1(n7205), .B2(n10167), .B3(n5728), .A(images_bus[418]), 
        .ZN(n10164) );
  aor22d1 U6232 ( .A1(n10387), .A2(n10388), .B1(n7370), .B2(n10169), .Z(n10155) );
  aoi31d1 U6235 ( .B1(images_bus[408]), .B2(n10151), .B3(images_bus[409]), .A(
        n12136), .ZN(n10157) );
  oai211d1 U6238 ( .C1(n5034), .C2(n10146), .A(images_bus[404]), .B(
        images_bus[405]), .ZN(n10149) );
  aon211d1 U6239 ( .C1(n10141), .C2(images_bus[399]), .B(n10389), .A(
        images_bus[402]), .ZN(n10146) );
  aoim21d1 U6240 ( .B1(n10137), .B2(n10135), .A(n6291), .ZN(n10141) );
  aoi21d1 U6244 ( .B1(n9447), .B2(n3221), .A(n7250), .ZN(n9604) );
  oan211d1 U6245 ( .C1(n6993), .C2(n8653), .B(n3233), .A(n6406), .ZN(n7250) );
  oai21d1 U6250 ( .B1(n3205), .B2(n10389), .A(n3193), .ZN(n8642) );
  aoi31d1 U6251 ( .B1(images_bus[393]), .B2(n10127), .B3(images_bus[392]), .A(
        n6837), .ZN(n10131) );
  aoim31d1 U6254 ( .B1(n10390), .B2(n12139), .B3(n4649), .A(n6366), .ZN(n10123) );
  oai21d1 U6255 ( .B1(n10390), .B2(n8621), .A(n10391), .ZN(n10121) );
  oai21d1 U6256 ( .B1(n10392), .B2(n12124), .A(n8621), .ZN(n10391) );
  oai31d1 U6268 ( .B1(n7154), .B2(images_bus[358]), .B3(n7161), .A(n6908), 
        .ZN(n10087) );
  aoi211d1 U6274 ( .C1(images_bus[323]), .C2(n10056), .A(n6606), .B(n4663), 
        .ZN(n10058) );
  aoi21d1 U6276 ( .B1(n3333), .B2(n9613), .A(n6919), .ZN(n10056) );
  aor31d1 U6280 ( .B1(images_bus[317]), .B2(n10040), .B3(images_bus[316]), .A(
        n6170), .Z(n10047) );
  oai31d1 U6284 ( .B1(n5405), .B2(n10038), .B3(n7006), .A(images_bus[314]), 
        .ZN(n10041) );
  aoi211d1 U6287 ( .C1(images_bus[307]), .C2(n10031), .A(n12146), .B(n4307), 
        .ZN(n10394) );
  aoim31d1 U6289 ( .B1(n5531), .B2(n10029), .B3(n7072), .A(n6752), .ZN(n10031)
         );
  aoi31d1 U6291 ( .B1(images_bus[300]), .B2(n3483), .B3(images_bus[301]), .A(
        n6303), .ZN(n10030) );
  aoim31d1 U6300 ( .B1(n7237), .B2(n10007), .B3(n5738), .A(n12122), .ZN(n10014) );
  oai211d1 U6307 ( .C1(n12169), .C2(n10001), .A(n6466), .B(images_bus[285]), 
        .ZN(n10004) );
  oai31d1 U6308 ( .B1(n5410), .B2(n10395), .B3(n7016), .A(images_bus[282]), 
        .ZN(n10001) );
  aon211d1 U6311 ( .C1(n9999), .C2(images_bus[275]), .B(n10397), .A(
        images_bus[278]), .ZN(n10396) );
  aoi31d1 U6312 ( .B1(images_bus[273]), .B2(n3507), .B3(images_bus[272]), .A(
        n6753), .ZN(n9999) );
  aoi311d1 U6314 ( .C1(images_bus[268]), .C2(n9986), .C3(images_bus[269]), .A(
        n6305), .B(n5933), .ZN(n9990) );
  aon211d1 U6316 ( .C1(n9980), .C2(images_bus[263]), .B(n9982), .A(
        images_bus[266]), .ZN(n9987) );
  oan211d1 U6317 ( .C1(n10398), .C2(n5266), .B(n9621), .A(n6388), .ZN(n9980)
         );
  aon211d1 U6321 ( .C1(n10403), .C2(n10398), .B(n6113), .A(n5348), .ZN(n9971)
         );
  aon211d1 U6322 ( .C1(n10404), .C2(images_bus[255]), .B(n10405), .A(
        images_bus[258]), .ZN(n10398) );
  aoi211d1 U6324 ( .C1(images_bus[251]), .C2(n9967), .A(n6469), .B(n3577), 
        .ZN(n9968) );
  aoi31d1 U6325 ( .B1(images_bus[249]), .B2(n9964), .B3(images_bus[248]), .A(
        n6677), .ZN(n9967) );
  aoi31d1 U6328 ( .B1(images_bus[245]), .B2(n9960), .B3(images_bus[244]), .A(
        n6246), .ZN(n9963) );
  aon211d1 U6329 ( .C1(n3799), .C2(n9960), .B(n6759), .A(n10407), .ZN(n9955)
         );
  oai311d1 U6330 ( .C1(n7076), .C2(n9951), .C3(n5542), .A(images_bus[243]), 
        .B(images_bus[242]), .ZN(n9960) );
  aoi211d1 U6333 ( .C1(images_bus[235]), .C2(n9944), .A(n4451), .B(n6567), 
        .ZN(n10408) );
  aoi21d1 U6335 ( .B1(n9941), .B2(n5652), .A(n6855), .ZN(n9944) );
  oai211d1 U6340 ( .C1(n5268), .C2(n9936), .A(n6621), .B(images_bus[229]), 
        .ZN(n9946) );
  oai31d1 U6341 ( .B1(n5747), .B2(n9934), .B3(n7242), .A(n6931), .ZN(n9936) );
  oai31d1 U6343 ( .B1(n3619), .B2(n9928), .B3(n6475), .A(images_bus[222]), 
        .ZN(n9931) );
  aoi31d1 U6345 ( .B1(images_bus[216]), .B2(n9923), .B3(images_bus[217]), .A(
        n12134), .ZN(n9930) );
  oai211d1 U6347 ( .C1(n5068), .C2(n9918), .A(images_bus[212]), .B(
        images_bus[213]), .ZN(n9921) );
  aoim31d1 U6352 ( .B1(n4459), .B2(n9907), .B3(n6571), .A(n12155), .ZN(n9913)
         );
  aoi311d1 U6355 ( .C1(images_bus[200]), .C2(n9904), .C3(images_bus[201]), .A(
        n12128), .B(n5186), .ZN(n9907) );
  oai21d1 U6357 ( .B1(n5276), .B2(n3812), .A(n7420), .ZN(n9901) );
  aoi21d1 U6360 ( .B1(n9894), .B2(n5756), .A(n6934), .ZN(n9895) );
  aoim31d1 U6363 ( .B1(n3814), .B2(n9887), .B3(n6481), .A(n12159), .ZN(n9891)
         );
  oai21d1 U6365 ( .B1(n9884), .B2(n9886), .A(images_bus[186]), .ZN(n9889) );
  aoi211d1 U6368 ( .C1(images_bus[179]), .C2(n9880), .A(n12145), .B(n4316), 
        .ZN(n9883) );
  aoi211d1 U6370 ( .C1(images_bus[175]), .C2(n9870), .A(n7081), .B(n5558), 
        .ZN(n10411) );
  aoi31d1 U6373 ( .B1(images_bus[173]), .B2(n9868), .B3(images_bus[172]), .A(
        n12154), .ZN(n9870) );
  or02d0 U6376 ( .A1(n9863), .A2(n6039), .Z(n9862) );
  oai21d1 U6378 ( .B1(n9859), .B2(n10412), .A(images_bus[166]), .ZN(n9863) );
  oai21d1 U6381 ( .B1(n9850), .B2(n10413), .A(images_bus[162]), .ZN(n9855) );
  aoi211d1 U6384 ( .C1(n9842), .C2(n9846), .A(n6484), .B(n3903), .ZN(n9853) );
  aoim31d1 U6389 ( .B1(n4319), .B2(n12144), .B3(n9835), .A(n6264), .ZN(n9840)
         );
  oai31d1 U6395 ( .B1(n7093), .B2(n9830), .B3(n5573), .A(images_bus[146]), 
        .ZN(n9834) );
  aoi211d1 U6398 ( .C1(images_bus[139]), .C2(n9823), .A(n6575), .B(n4491), 
        .ZN(n10415) );
  aoi31d1 U6399 ( .B1(images_bus[137]), .B2(n9826), .B3(images_bus[136]), .A(
        n12127), .ZN(n9823) );
  oai21d1 U6401 ( .B1(n9817), .B2(n10416), .A(images_bus[134]), .ZN(n9827) );
  aoi211d1 U6402 ( .C1(n3985), .C2(n5771), .A(n6946), .B(n5281), .ZN(n9817) );
  aoi211d1 U6407 ( .C1(images_bus[123]), .C2(n9812), .A(n6488), .B(n3986), 
        .ZN(n9815) );
  oai211d1 U6409 ( .C1(n5855), .C2(n4059), .A(images_bus[120]), .B(
        images_bus[121]), .ZN(n10417) );
  oan211d1 U6411 ( .C1(n9801), .C2(n5104), .B(n9072), .A(n6267), .ZN(n9807) );
  oai211d1 U6413 ( .C1(n5957), .C2(n9797), .A(images_bus[112]), .B(
        images_bus[113]), .ZN(n10418) );
  oai211d1 U6415 ( .C1(n5203), .C2(n4060), .A(images_bus[109]), .B(
        images_bus[108]), .ZN(n10419) );
  aoi31d1 U6417 ( .B1(images_bus[105]), .B2(n9786), .B3(images_bus[104]), .A(
        n6875), .ZN(n9790) );
  oaim22d1 U6422 ( .A1(images_bus[102]), .A2(n9050), .B1(n9786), .B2(n6787), 
        .ZN(n9781) );
  oai211d1 U6424 ( .C1(n5284), .C2(n9782), .A(images_bus[100]), .B(
        images_bus[101]), .ZN(n10420) );
  nd13d1 U6426 ( .A1(n9779), .A2(images_bus[96]), .A3(images_bus[97]), .ZN(
        n9785) );
  aoi211d1 U6428 ( .C1(images_bus[91]), .C2(n9767), .A(n12148), .B(n4119), 
        .ZN(n9775) );
  oai211d1 U6431 ( .C1(n5858), .C2(n9763), .A(images_bus[88]), .B(
        images_bus[89]), .ZN(n10421) );
  oai211d1 U6433 ( .C1(n5106), .C2(n9764), .A(images_bus[84]), .B(
        images_bus[85]), .ZN(n10422) );
  oai31d1 U6434 ( .B1(n5581), .B2(n9758), .B3(n7104), .A(images_bus[82]), .ZN(
        n9764) );
  oai31d1 U6436 ( .B1(n6586), .B2(n9753), .B3(n4503), .A(images_bus[78]), .ZN(
        n9757) );
  aoi31d1 U6441 ( .B1(images_bus[69]), .B2(n9745), .B3(images_bus[68]), .A(
        n6403), .ZN(n9748) );
  aoim21d1 U6444 ( .B1(n9738), .B2(n5803), .A(n6953), .ZN(n9743) );
  aor31d1 U6448 ( .B1(images_bus[60]), .B2(n9732), .B3(images_bus[61]), .A(
        n6200), .Z(n9735) );
  oai211d1 U6450 ( .C1(n5862), .C2(n9720), .A(images_bus[56]), .B(
        images_bus[57]), .ZN(n9729) );
  oai31d1 U6453 ( .B1(n6550), .B2(n12172), .B3(n9719), .A(images_bus[54]), 
        .ZN(n9720) );
  aoim31d1 U6456 ( .B1(n5585), .B2(n9713), .B3(n7105), .A(n12130), .ZN(n9715)
         );
  oai211d1 U6460 ( .C1(n6070), .C2(n9703), .A(images_bus[40]), .B(
        images_bus[41]), .ZN(n9706) );
  or02d0 U6461 ( .A1(n10425), .A2(n6411), .Z(n9703) );
  aoi211d1 U6462 ( .C1(images_bus[35]), .C2(n9701), .A(n6646), .B(n4754), .ZN(
        n10425) );
  aoi21d1 U6463 ( .B1(n9695), .B2(n5784), .A(n12120), .ZN(n9701) );
  nd13d1 U6465 ( .A1(n9690), .A2(images_bus[30]), .A3(images_bus[31]), .ZN(
        n9695) );
  aoi211d1 U6466 ( .C1(images_bus[27]), .C2(n4347), .A(n6507), .B(n4292), .ZN(
        n9690) );
  oai211d1 U6472 ( .C1(n5864), .C2(n4352), .A(images_bus[25]), .B(
        images_bus[24]), .ZN(n10427) );
  aoi31d1 U6475 ( .B1(images_bus[20]), .B2(n10428), .B3(images_bus[21]), .A(
        n6273), .ZN(n9677) );
  oai211d1 U6477 ( .C1(n5591), .C2(n10429), .A(images_bus[19]), .B(
        images_bus[18]), .ZN(n10428) );
  aor31d1 U6478 ( .B1(images_bus[15]), .B2(n9665), .B3(images_bus[14]), .A(
        n7109), .Z(n10429) );
  oai211d1 U6480 ( .C1(n5220), .C2(n9660), .A(images_bus[12]), .B(
        images_bus[13]), .ZN(n9665) );
  aon211d1 U6481 ( .C1(n9649), .C2(images_bus[7]), .B(n8903), .A(n6890), .ZN(
        n9660) );
  oan211d1 U6483 ( .C1(n5315), .C2(n6975), .B(n8897), .A(n6413), .ZN(n9649) );
  oai21d1 U6487 ( .B1(images_bus[1]), .B2(n5008), .A(n10432), .ZN(N26358) );
  oan211d1 U6489 ( .C1(n10434), .C2(n9652), .B(n10435), .A(n5785), .ZN(n10433)
         );
  aoi22d1 U6490 ( .A1(n4854), .A2(n10436), .B1(n8894), .B2(n10437), .ZN(n10434) );
  oai311d1 U6491 ( .C1(n4771), .C2(n10438), .C3(n9661), .A(n9656), .B(n10439), 
        .ZN(n10436) );
  aoi22d1 U6492 ( .A1(n4766), .A2(n10440), .B1(images_bus[6]), .B2(n10437), 
        .ZN(n10439) );
  aoi31d1 U6494 ( .B1(N8107), .B2(n10442), .B3(n4816), .A(n4881), .ZN(n10438)
         );
  oai22d1 U6495 ( .A1(n10444), .A2(n10445), .B1(n10446), .B2(n10430), .ZN(
        n10442) );
  aoi311d1 U6496 ( .C1(n4604), .C2(n10447), .C3(n4628), .A(n4608), .B(n10448), 
        .ZN(n10446) );
  aoi311d1 U6497 ( .C1(n10449), .C2(n10450), .C3(n10451), .A(n7462), .B(n10452), .ZN(n10448) );
  aon211d1 U6500 ( .C1(n4568), .C2(n10455), .B(n10456), .A(n7472), .ZN(n10451)
         );
  oan211d1 U6501 ( .C1(n4549), .C2(n6552), .B(n10458), .A(n10459), .ZN(n10456)
         );
  aoim31d1 U6502 ( .B1(n7485), .B2(n4361), .B3(n10460), .A(n10461), .ZN(n10458) );
  oan211d1 U6503 ( .C1(n10462), .C2(n9679), .B(images_bus[21]), .A(n10463), 
        .ZN(n10461) );
  aon211d1 U6504 ( .C1(n8161), .C2(n10464), .B(n10465), .A(n4576), .ZN(n10460)
         );
  aoi311d1 U6505 ( .C1(n10466), .C2(n10467), .C3(images_bus[27]), .A(n9687), 
        .B(n9684), .ZN(n10465) );
  aon211d1 U6506 ( .C1(n10468), .C2(n10469), .B(n10470), .A(n4376), .ZN(n10466) );
  aoi221d1 U6508 ( .B1(n4281), .B2(n6146), .C1(n4278), .C2(n10475), .A(n10476), 
        .ZN(n10471) );
  oai22d1 U6509 ( .A1(n10477), .A2(n10478), .B1(n10479), .B2(n4231), .ZN(
        n10475) );
  aoi311d1 U6510 ( .C1(n6691), .C2(n10480), .C3(n10481), .A(n10482), .B(n4243), 
        .ZN(n10479) );
  oaim22d1 U6511 ( .A1(n12120), .A2(n10477), .B1(n10484), .B2(n4233), .ZN(
        n10482) );
  aoi21d1 U6512 ( .B1(images_bus[39]), .B2(n10485), .A(n10486), .ZN(n10481) );
  oai211d1 U6513 ( .C1(n10487), .C2(n10488), .A(n10489), .B(n4274), .ZN(n10485) );
  oan211d1 U6515 ( .C1(n10490), .C2(n10491), .B(n10492), .A(n10493), .ZN(
        n10487) );
  aoi221d1 U6516 ( .B1(images_bus[44]), .B2(n4295), .C1(n4249), .C2(n10496), 
        .A(n8950), .ZN(n10490) );
  oaim22d1 U6519 ( .A1(n10497), .A2(n9714), .B1(n10498), .B2(n4271), .ZN(
        n10496) );
  aoi31d1 U6520 ( .B1(n6720), .B2(n10499), .B3(n7511), .A(n6724), .ZN(n10497)
         );
  oai31d1 U6521 ( .B1(n10500), .B2(n10501), .B3(n5110), .A(n4294), .ZN(n10499)
         );
  aoi311d1 U6522 ( .C1(n8216), .C2(n10503), .C3(n4259), .A(n10504), .B(n10505), 
        .ZN(n10501) );
  aoi311d1 U6523 ( .C1(n10506), .C2(n10507), .C3(images_bus[55]), .A(n8974), 
        .B(n10508), .ZN(n10505) );
  aon211d1 U6524 ( .C1(n4262), .C2(n10509), .B(n10510), .A(n9726), .ZN(n10506)
         );
  aoim21d1 U6525 ( .B1(n10511), .B2(n10512), .A(n6730), .ZN(n10510) );
  oai22d1 U6526 ( .A1(n4293), .A2(n6701), .B1(n10514), .B2(n8116), .ZN(n10512)
         );
  oai211d1 U6527 ( .C1(n10515), .C2(n5799), .A(n10516), .B(n8227), .ZN(n10511)
         );
  oai211d1 U6529 ( .C1(n10520), .C2(n5810), .A(n10521), .B(images_bus[67]), 
        .ZN(n10519) );
  aoim211d1 U6531 ( .C1(n9004), .C2(n10522), .A(n10523), .B(n10524), .ZN(
        n10520) );
  aon211d1 U6532 ( .C1(n10525), .C2(n10526), .B(n10527), .A(n10528), .ZN(
        n10523) );
  aon211d1 U6536 ( .C1(images_bus[76]), .C2(n10530), .B(n10532), .A(n4151), 
        .ZN(n10526) );
  oai21d1 U6540 ( .B1(n4155), .B2(n10533), .A(n4156), .ZN(n10532) );
  aon211d1 U6542 ( .C1(n10534), .C2(n4179), .B(n10535), .A(n4178), .ZN(n10533)
         );
  oan211d1 U6543 ( .C1(n10536), .C2(n10537), .B(n4140), .A(n5958), .ZN(n10534)
         );
  aoi321d1 U6544 ( .C1(n4159), .C2(n4163), .C3(n10540), .B1(n4176), .B2(n10541), .A(n5842), .ZN(n10536) );
  oai22d1 U6546 ( .A1(n10543), .A2(n10544), .B1(n10545), .B2(n4158), .ZN(
        n10541) );
  oan211d1 U6548 ( .C1(n10546), .C2(n5859), .B(n10547), .A(n6268), .ZN(n10540)
         );
  oan211d1 U6549 ( .C1(n8881), .C2(n10548), .B(n8266), .A(n10549), .ZN(n10547)
         );
  oan211d1 U6550 ( .C1(n4120), .C2(n5027), .B(n10551), .A(n5037), .ZN(n10549)
         );
  aon211d1 U6553 ( .C1(n4117), .C2(n10552), .B(n10553), .A(n8105), .ZN(n10551)
         );
  oai321d1 U6554 ( .C1(n5882), .C2(n10554), .C3(n10555), .B1(n10556), .B2(
        n5031), .A(n10557), .ZN(n10552) );
  aoim31d1 U6555 ( .B1(n10558), .B2(n6786), .B3(n5019), .A(n10559), .ZN(n10556) );
  aoi221d1 U6557 ( .B1(n4068), .B2(n10560), .C1(n6787), .C2(n10561), .A(n4745), 
        .ZN(n10558) );
  oai321d1 U6558 ( .C1(n9791), .C2(n10562), .C3(n7578), .B1(images_bus[105]), 
        .B2(n5905), .A(n10563), .ZN(n10560) );
  aoi31d1 U6559 ( .B1(n5911), .B2(n10564), .B3(n4072), .A(n10565), .ZN(n10563)
         );
  oai22d1 U6564 ( .A1(n10566), .A2(n5915), .B1(n10567), .B2(n9795), .ZN(n10564) );
  aoi321d1 U6566 ( .C1(n10568), .C2(n10569), .C3(n4081), .B1(n4104), .B2(
        n10571), .A(n10572), .ZN(n10567) );
  oai311d1 U6570 ( .C1(n7590), .C2(n4121), .C3(n9071), .A(n9799), .B(n10574), 
        .ZN(n10569) );
  aoi22d1 U6571 ( .A1(n5036), .A2(n10575), .B1(n10571), .B2(n6795), .ZN(n10574) );
  oai211d1 U6572 ( .C1(n4121), .C2(n6267), .A(n10576), .B(n7439), .ZN(n10575)
         );
  aon211d1 U6573 ( .C1(n10577), .C2(n4093), .B(n10579), .A(n9073), .ZN(n10576)
         );
  oan211d1 U6575 ( .C1(n10580), .C2(n6829), .B(n10581), .A(n5447), .ZN(n10577)
         );
  oai211d1 U6576 ( .C1(n10582), .C2(n10583), .A(n4092), .B(n4096), .ZN(n10581)
         );
  oan211d1 U6579 ( .C1(n10585), .C2(n4002), .B(n10586), .A(n5041), .ZN(n10582)
         );
  aoi221d1 U6584 ( .B1(n4391), .B2(n10588), .C1(n4004), .C2(n3988), .A(n10590), 
        .ZN(n10585) );
  oai222d1 U6585 ( .A1(images_bus[133]), .A2(n9638), .B1(n10591), .B2(n5055), 
        .C1(n10592), .C2(n6848), .ZN(n10588) );
  oan211d1 U6592 ( .C1(n10594), .C2(n10595), .B(n6851), .A(n10595), .ZN(n10591) );
  oan211d1 U6593 ( .C1(n10596), .C2(n8321), .B(n10597), .A(n6853), .ZN(n10594)
         );
  oai31d1 U6594 ( .B1(n10598), .B2(n10599), .B3(n10600), .A(n4017), .ZN(n10597) );
  aoi311d1 U6597 ( .C1(n10604), .C2(n10605), .C3(n10606), .A(n4023), .B(n6860), 
        .ZN(n10600) );
  aoi21d1 U6600 ( .B1(n5081), .B2(n10607), .A(n10608), .ZN(n10606) );
  aon211d1 U6602 ( .C1(n4048), .C2(n10610), .B(n10611), .A(n4028), .ZN(n10605)
         );
  oai22d1 U6607 ( .A1(n10615), .A2(n4389), .B1(n10616), .B2(n7437), .ZN(n10610) );
  aoi221d1 U6612 ( .B1(n6868), .B2(n10618), .C1(n4039), .C2(n10619), .A(n10620), .ZN(n10616) );
  oai211d1 U6613 ( .C1(n10621), .C2(n4418), .A(n10622), .B(n10623), .ZN(n10618) );
  aoi22d1 U6614 ( .A1(n3909), .A2(n10624), .B1(images_bus[156]), .B2(n10619), 
        .ZN(n10623) );
  aoi31d1 U6615 ( .B1(n5120), .B2(n5762), .B3(n3908), .A(n9122), .ZN(n10622)
         );
  aoi22d1 U6626 ( .A1(n10627), .A2(n6883), .B1(n3914), .B2(n10628), .ZN(n10621) );
  oan211d1 U6628 ( .C1(n10629), .C2(n10630), .B(n10631), .A(n10632), .ZN(
        n10627) );
  aoi31d1 U6629 ( .B1(n3920), .B2(n10633), .B3(n3922), .A(n10634), .ZN(n10631)
         );
  oan211d1 U6630 ( .C1(n10635), .C2(n5144), .B(n10636), .A(n5132), .ZN(n10634)
         );
  oai322d1 U6632 ( .C1(n6899), .C2(n3904), .C3(n10640), .A1(n10641), .A2(n9872), .B1(n10642), .B2(n10643), .ZN(n10638) );
  aoi311d1 U6636 ( .C1(n6910), .C2(n10644), .C3(n9632), .A(n10645), .B(n9875), 
        .ZN(n10641) );
  oai22d1 U6637 ( .A1(n12154), .A2(n3904), .B1(n3905), .B2(n5158), .ZN(n10645)
         );
  oai221d1 U6640 ( .B1(n3905), .B2(n10648), .C1(n10649), .C2(n5999), .A(n9879), 
        .ZN(n10644) );
  aoi211d1 U6643 ( .C1(n6003), .C2(n10650), .A(n10651), .B(n10652), .ZN(n10649) );
  aoi311d1 U6644 ( .C1(n10653), .C2(n10654), .C3(n10655), .A(n5177), .B(n3954), 
        .ZN(n10652) );
  aoi31d1 U6647 ( .B1(n8383), .B2(n10658), .B3(n9144), .A(n10659), .ZN(n10655)
         );
  oai222d1 U6651 ( .A1(n3906), .A2(n6481), .B1(n10662), .B2(n10663), .C1(n3828), .C2(n5187), .ZN(n10658) );
  oan211d1 U6652 ( .C1(n10664), .C2(n10665), .B(n3820), .A(n10667), .ZN(n10662) );
  oaim21d1 U6655 ( .B1(n6179), .B2(n10667), .A(images_bus[191]), .ZN(n10665)
         );
  oai322d1 U6656 ( .C1(n10668), .C2(n3837), .C3(n8391), .A1(n10669), .A2(n4390), .B1(n3815), .B2(n6014), .ZN(n10664) );
  aoi321d1 U6658 ( .C1(n3836), .C2(n6038), .C3(n3833), .B1(n3834), .B2(n10673), 
        .A(n5276), .ZN(n10669) );
  aon211d1 U6665 ( .C1(n3844), .C2(n10677), .B(n10678), .A(n3822), .ZN(n10668)
         );
  oai221d1 U6671 ( .B1(n10679), .B2(n10680), .C1(n12128), .C2(n3816), .A(
        n10682), .ZN(n10677) );
  oan211d1 U6673 ( .C1(n10686), .C2(n4388), .B(n10687), .A(n10688), .ZN(n10684) );
  or02d0 U6674 ( .A1(n5225), .A2(n6951), .Z(n4388) );
  aoi311d1 U6675 ( .C1(n5232), .C2(n10689), .C3(n3875), .A(n10690), .B(n10691), 
        .ZN(n10686) );
  aoi221d1 U6679 ( .B1(n3856), .B2(n10694), .C1(n3872), .C2(n10696), .A(n10689), .ZN(n10692) );
  oai22d1 U6680 ( .A1(n10697), .A2(n7418), .B1(n10698), .B2(n8416), .ZN(n10694) );
  aoim211d1 U6681 ( .C1(n7019), .C2(n10697), .A(n3860), .B(n10699), .ZN(n10698) );
  oan211d1 U6682 ( .C1(n10700), .C2(n10701), .B(n10702), .A(n8423), .ZN(n10699) );
  aon211d1 U6684 ( .C1(n9189), .C2(n10703), .B(n10704), .A(n3864), .ZN(n10701)
         );
  oai321d1 U6685 ( .C1(n3730), .C2(n10706), .C3(n10707), .B1(n3664), .B2(n3732), .A(n10710), .ZN(n10703) );
  aoi221d1 U6686 ( .B1(n10711), .B2(n6931), .C1(n3742), .C2(n5268), .A(n10712), 
        .ZN(n10706) );
  oai322d1 U6687 ( .C1(n9940), .C2(n10713), .C3(n9202), .A1(n10714), .A2(n4401), .B1(n10715), .B2(n9194), .ZN(n10712) );
  aoi22d1 U6691 ( .A1(n10716), .A2(n10717), .B1(n3761), .B2(n10718), .ZN(
        n10714) );
  aoi31d1 U6692 ( .B1(n10719), .B2(n10720), .B3(n10721), .A(n10722), .ZN(
        n10717) );
  aoi21d1 U6693 ( .B1(n8440), .B2(n10723), .A(n5173), .ZN(n10721) );
  aon211d1 U6695 ( .C1(n3801), .C2(n10724), .B(n10725), .A(n4420), .ZN(n10719)
         );
  aoi311d1 U6700 ( .C1(n3799), .C2(n3660), .C3(n9624), .A(n10730), .B(n10731), 
        .ZN(n10727) );
  oai22d1 U6701 ( .A1(images_bus[241]), .A2(n10732), .B1(n2811), .B2(n4417), 
        .ZN(n10730) );
  oai321d1 U6705 ( .C1(n9227), .C2(n10737), .C3(n7002), .B1(n6538), .B2(n10738), .A(n7004), .ZN(n10736) );
  aoim31d1 U6706 ( .B1(n5835), .B2(n10739), .B3(n5326), .A(n10740), .ZN(n10737) );
  aoi311d1 U6707 ( .C1(n3780), .C2(n10742), .C3(n3785), .A(n10740), .B(n10744), 
        .ZN(n10739) );
  aoi321d1 U6709 ( .C1(n3574), .C2(images_bus[254]), .C3(n10747), .B1(n3788), 
        .B2(n10748), .A(n3659), .ZN(n10745) );
  aoi31d1 U6711 ( .B1(n10751), .B2(n10752), .B3(n10753), .A(n3522), .ZN(n10747) );
  aoi22d1 U6712 ( .A1(n3525), .A2(n10755), .B1(n5348), .B2(n6113), .ZN(n10753)
         );
  oai211d1 U6713 ( .C1(n10756), .C2(n9243), .A(n10757), .B(n10758), .ZN(n10755) );
  aoim31d1 U6714 ( .B1(n3530), .B2(n10759), .B3(n9239), .A(n10760), .ZN(n10758) );
  or02d0 U6717 ( .A1(n10762), .A2(n10764), .Z(n8468) );
  aoi321d1 U6721 ( .C1(n7754), .C2(n10765), .C3(n8471), .B1(n5744), .B2(n10766), .A(n10767), .ZN(n10756) );
  aoi211d1 U6722 ( .C1(images_bus[265]), .C2(n10768), .A(n9981), .B(n3567), 
        .ZN(n10767) );
  oai211d1 U6723 ( .C1(n10770), .C2(n4456), .A(n10771), .B(n10772), .ZN(n10766) );
  aoi31d1 U6724 ( .B1(n10773), .B2(n10774), .B3(n3566), .A(n10775), .ZN(n10772) );
  aoi22d1 U6726 ( .A1(n3559), .A2(n10778), .B1(n10779), .B2(n10780), .ZN(
        n10776) );
  oaim22d1 U6727 ( .A1(n10781), .A2(n5359), .B1(n5359), .B2(n10779), .ZN(
        n10778) );
  oan211d1 U6728 ( .C1(n10782), .C2(n10783), .B(n3544), .A(n10785), .ZN(n10781) );
  oai22d1 U6732 ( .A1(n10788), .A2(n3582), .B1(n9617), .B2(n10790), .ZN(n10783) );
  oai211d1 U6734 ( .C1(images_bus[281]), .C2(n9617), .A(n10792), .B(n10793), 
        .ZN(n10782) );
  oai22d1 U6738 ( .A1(n10800), .A2(n8502), .B1(n3554), .B2(n10801), .ZN(n10799) );
  aoi321d1 U6739 ( .C1(n9273), .C2(n10794), .C3(images_bus[286]), .B1(n10802), 
        .B2(n3424), .A(n10803), .ZN(n10800) );
  oan211d1 U6741 ( .C1(n10805), .C2(n3475), .B(n10807), .A(n5382), .ZN(n10802)
         );
  aoi31d1 U6742 ( .B1(n3475), .B2(n10808), .B3(n8509), .A(n10809), .ZN(n10807)
         );
  oan211d1 U6743 ( .C1(n10805), .C2(n3474), .B(n10810), .A(n8510), .ZN(n10809)
         );
  oai321d1 U6748 ( .C1(n4495), .C2(n10813), .C3(n8507), .B1(n3471), .B2(n10814), .A(n10815), .ZN(n10808) );
  aoi311d1 U6750 ( .C1(n5396), .C2(n10816), .C3(images_bus[296]), .A(n10817), 
        .B(n10818), .ZN(n10813) );
  aon211d1 U6752 ( .C1(n10820), .C2(n10821), .B(n7783), .A(n10822), .ZN(n10817) );
  aoim31d1 U6760 ( .B1(n3439), .B2(n10827), .B3(n5404), .A(n8523), .ZN(n10821)
         );
  aoi22d1 U6763 ( .A1(n3432), .A2(n10829), .B1(n10830), .B2(n7078), .ZN(n10820) );
  oai322d1 U6764 ( .C1(n6181), .C2(n3436), .C3(n10831), .A1(n10832), .A2(n9303), .B1(n10827), .B2(n3438), .ZN(n10829) );
  aoi22d1 U6766 ( .A1(n10833), .A2(n3456), .B1(n7090), .B2(n10834), .ZN(n10832) );
  oan211d1 U6767 ( .C1(n3454), .C2(n10835), .B(n10836), .A(n7090), .ZN(n10833)
         );
  oai22d1 U6769 ( .A1(n10839), .A2(n9309), .B1(n10840), .B2(n10841), .ZN(
        n10838) );
  oai21d1 U6770 ( .B1(images_bus[312]), .B2(n9312), .A(n3450), .ZN(n10841) );
  aoi321d1 U6771 ( .C1(n10843), .C2(n9315), .C3(n10844), .B1(n10039), .B2(
        n10845), .A(n5826), .ZN(n10839) );
  oai322d1 U6773 ( .C1(n6675), .C2(n3443), .C3(n3485), .A1(n10847), .A2(n10848), .B1(n5418), .B2(n10849), .ZN(n10845) );
  aon211d1 U6774 ( .C1(n10850), .C2(n10851), .B(n10852), .A(n6194), .ZN(n10849) );
  aoi21d1 U6775 ( .B1(images_bus[319]), .B2(n10853), .A(n3360), .ZN(n10852) );
  aon211d1 U6778 ( .C1(n3366), .C2(n10855), .B(n10856), .A(n3363), .ZN(n10853)
         );
  oan211d1 U6782 ( .C1(n3418), .C2(n6919), .B(n3366), .A(n10859), .ZN(n10856)
         );
  oai322d1 U6783 ( .C1(n6203), .C2(n10860), .C3(n10861), .A1(n8549), .A2(
        n10862), .B1(images_bus[325]), .B2(n7817), .ZN(n10855) );
  aon211d1 U6786 ( .C1(images_bus[324]), .C2(n10863), .B(n4538), .A(n10864), 
        .ZN(n10862) );
  aoi31d1 U6787 ( .B1(n3410), .B2(n3372), .B3(n10866), .A(n10867), .ZN(n10860)
         );
  aoi211d1 U6789 ( .C1(images_bus[329]), .C2(n10870), .A(n10869), .B(n10863), 
        .ZN(n10866) );
  aon211d1 U6790 ( .C1(n3405), .C2(n10871), .B(n10872), .A(n3409), .ZN(n10870)
         );
  oai311d1 U6792 ( .C1(n10874), .C2(n10875), .C3(n3378), .A(n10876), .B(n10877), .ZN(n10871) );
  aoi31d1 U6793 ( .B1(n3376), .B2(n10879), .B3(n3374), .A(n10880), .ZN(n10877)
         );
  aoi322d1 U6799 ( .C1(images_bus[338]), .C2(n10879), .C3(n10886), .A1(n7135), 
        .A2(n10887), .B1(n3399), .B2(n5046), .ZN(n10875) );
  oai211d1 U6800 ( .C1(n10888), .C2(n7141), .A(n10889), .B(n10890), .ZN(n10887) );
  aoi22d1 U6801 ( .A1(n3334), .A2(n10892), .B1(n10893), .B2(n6258), .ZN(n10890) );
  aon211d1 U6802 ( .C1(n3396), .C2(n5825), .B(n3334), .A(n10895), .ZN(n10889)
         );
  oai21d1 U6803 ( .B1(n3393), .B2(n6998), .A(n3395), .ZN(n10895) );
  aoi31d1 U6808 ( .B1(n9363), .B2(n10898), .B3(n3393), .A(n10899), .ZN(n10888)
         );
  oan211d1 U6809 ( .C1(n8570), .C2(n10900), .B(n10901), .A(n7139), .ZN(n10899)
         );
  oan211d1 U6810 ( .C1(n10902), .C2(n10903), .B(n7142), .A(n10904), .ZN(n10901) );
  aon211d1 U6812 ( .C1(images_bus[350]), .C2(n10086), .B(n6281), .A(n10906), 
        .ZN(n10905) );
  oan211d1 U6814 ( .C1(n3330), .C2(n7222), .B(n3273), .A(n10907), .ZN(n10903)
         );
  aoi22d1 U6816 ( .A1(n10911), .A2(n10912), .B1(n3275), .B2(n10913), .ZN(
        n10908) );
  oai22d1 U6817 ( .A1(n10914), .A2(n4586), .B1(n10915), .B2(n10090), .ZN(
        n10913) );
  aoi322d1 U6818 ( .C1(n5477), .C2(n6601), .C3(n10916), .A1(n3323), .A2(n4653), 
        .B1(n10917), .B2(n3320), .ZN(n10914) );
  oan211d1 U6819 ( .C1(n10918), .C2(n10919), .B(n10920), .A(n7857), .ZN(n10917) );
  aoi31d1 U6820 ( .B1(n3316), .B2(n10921), .B3(n5480), .A(n10922), .ZN(n10920)
         );
  oai211d1 U6823 ( .C1(n7381), .C2(n10925), .A(n10926), .B(n10927), .ZN(n10921) );
  aon211d1 U6824 ( .C1(n3286), .C2(n5920), .B(n10928), .A(n5486), .ZN(n10927)
         );
  oan211d1 U6828 ( .C1(n10929), .C2(n7180), .B(n10930), .A(n10931), .ZN(n10928) );
  oai211d1 U6829 ( .C1(images_bus[368]), .C2(n10932), .A(n10102), .B(n10933), 
        .ZN(n10930) );
  or02d0 U6832 ( .A1(n10102), .A2(n10097), .Z(n7180) );
  aoi22d1 U6834 ( .A1(n10936), .A2(n5491), .B1(n3291), .B2(n10937), .ZN(n10929) );
  aon211d1 U6835 ( .C1(n10938), .C2(n10939), .B(n5492), .A(n6327), .ZN(n10937)
         );
  aoi321d1 U6838 ( .C1(n10940), .C2(n10941), .C3(n10942), .B1(n3310), .B2(
        n10944), .A(n10945), .ZN(n10939) );
  aoi22d1 U6843 ( .A1(n5504), .A2(n3312), .B1(n5501), .B2(n10106), .ZN(n9398)
         );
  oai211d1 U6845 ( .C1(n10951), .C2(n10952), .A(n10106), .B(n10953), .ZN(n9404) );
  oai321d1 U6847 ( .C1(n6593), .C2(n10954), .C3(n10955), .B1(n10956), .B2(
        n9410), .A(n10957), .ZN(n10949) );
  aoi22d1 U6850 ( .A1(n3250), .A2(n10960), .B1(n6365), .B2(n10961), .ZN(n10956) );
  oai321d1 U6851 ( .C1(n8621), .C2(n10962), .C3(n10963), .B1(n3249), .B2(
        n10965), .A(n10966), .ZN(n10960) );
  aor211d1 U6852 ( .C1(n10965), .C2(images_bus[385]), .A(n7217), .B(n6364), 
        .Z(n10966) );
  aoi321d1 U6853 ( .C1(n10967), .C2(n7606), .C3(n10969), .B1(n9421), .B2(n4649), .A(n10970), .ZN(n10962) );
  oai22d1 U6854 ( .A1(n10969), .A2(n3137), .B1(n10972), .B2(n7223), .ZN(n10970) );
  aoi22d1 U6855 ( .A1(n10973), .A2(n3174), .B1(n6372), .B2(n10967), .ZN(n10972) );
  oan211d1 U6856 ( .C1(n10975), .C2(n3243), .B(n10976), .A(n8620), .ZN(n10973)
         );
  aoi31d1 U6857 ( .B1(n9425), .B2(n10977), .B3(n3243), .A(n10978), .ZN(n10976)
         );
  aoi221d1 U6859 ( .B1(n10980), .B2(n10138), .C1(n7230), .C2(n10981), .A(
        n10982), .ZN(n10979) );
  aon211d1 U6861 ( .C1(n3193), .C2(n3241), .B(n3135), .A(n10986), .ZN(n10981)
         );
  aoi31d1 U6862 ( .B1(n7235), .B2(n5906), .B3(n3241), .A(n10987), .ZN(n10986)
         );
  oan211d1 U6863 ( .C1(n10988), .C2(n3205), .B(n10989), .A(n7893), .ZN(n10987)
         );
  aoi22d1 U6865 ( .A1(n3204), .A2(n10990), .B1(n10991), .B2(n8836), .ZN(n10989) );
  aon211d1 U6866 ( .C1(images_bus[403]), .C2(n3136), .B(n8837), .A(n10993), 
        .ZN(n10990) );
  aon211d1 U6867 ( .C1(n3208), .C2(n10994), .B(n10995), .A(n3236), .ZN(n10993)
         );
  oan211d1 U6869 ( .C1(n3232), .C2(n6225), .B(n3208), .A(n10997), .ZN(n10995)
         );
  oai222d1 U6870 ( .A1(n10998), .A2(n10999), .B1(n3216), .B2(n11001), .C1(
        n11002), .C2(n8056), .ZN(n10994) );
  aoi221d1 U6872 ( .B1(n11004), .B2(n10388), .C1(n11005), .C2(n3226), .A(
        n11007), .ZN(n11002) );
  aoi22d1 U6874 ( .A1(n8682), .A2(n11011), .B1(n3038), .B2(n11012), .ZN(n11008) );
  oai321d1 U6875 ( .C1(n3046), .C2(n11013), .C3(n4713), .B1(n8672), .B2(n11014), .A(n11015), .ZN(n11012) );
  or04d0 U6876 ( .A1(n3042), .A2(n11016), .A3(n8683), .A4(n11017), .Z(n11015)
         );
  aon211d1 U6881 ( .C1(images_bus[418]), .C2(n6577), .B(n10386), .A(n11018), 
        .ZN(n11014) );
  aoi322d1 U6882 ( .C1(n3127), .C2(n3126), .C3(n11020), .A1(n11021), .A2(
        n11022), .B1(n4729), .B2(n11023), .ZN(n11013) );
  aoi31d1 U6883 ( .B1(n9464), .B2(N14242), .B3(n2812), .A(n11025), .ZN(n11020)
         );
  oan211d1 U6884 ( .C1(n5980), .C2(n11026), .B(N14242), .A(n11021), .ZN(n11025) );
  oai31d1 U6886 ( .B1(n9468), .B2(n11027), .B3(n8692), .A(n11028), .ZN(n11026)
         );
  aon211d1 U6887 ( .C1(n3064), .C2(n11029), .B(n11030), .A(n10181), .ZN(n11028) );
  aon211d1 U6889 ( .C1(n3062), .C2(n3123), .B(n11032), .A(n11033), .ZN(n11030)
         );
  oai21d1 U6892 ( .B1(n12142), .B2(n3069), .A(n3066), .ZN(n7952) );
  oai22d1 U6895 ( .A1(n11036), .A2(n5597), .B1(n11037), .B2(n11038), .ZN(
        n11029) );
  aon211d1 U6896 ( .C1(images_bus[430]), .C2(n10188), .B(n11039), .A(n11040), 
        .ZN(n11038) );
  aoi311d1 U6897 ( .C1(n3081), .C2(n3113), .C3(n11041), .A(n11042), .B(n11043), 
        .ZN(n11036) );
  oan211d1 U6898 ( .C1(n11044), .C2(n3083), .B(n11046), .A(n3119), .ZN(n11043)
         );
  aon211d1 U6901 ( .C1(images_bus[434]), .C2(n6564), .B(n9602), .A(n11048), 
        .ZN(n11046) );
  aoi321d1 U6905 ( .C1(n11049), .C2(n4300), .C3(n9599), .B1(n8716), .B2(n11050), .A(n11051), .ZN(n11044) );
  oai31d1 U6906 ( .B1(n11052), .B2(n6519), .B3(n11053), .A(n11054), .ZN(n11051) );
  oai21d1 U6908 ( .B1(n11056), .B2(n11049), .A(n3020), .ZN(n11052) );
  oai211d1 U6909 ( .C1(n3108), .C2(n11058), .A(n11059), .B(n11060), .ZN(n11050) );
  aon211d1 U6913 ( .C1(n7300), .C2(n11063), .B(n11064), .A(n3108), .ZN(n11059)
         );
  aon211d1 U6914 ( .C1(n11058), .C2(n5354), .B(n11065), .A(n11066), .ZN(n11064) );
  aon211d1 U6915 ( .C1(n11067), .C2(n6500), .B(n11068), .A(n5619), .ZN(n11066)
         );
  oan211d1 U6916 ( .C1(n3105), .C2(n6428), .B(n3103), .A(n3019), .ZN(n11068)
         );
  oan211d1 U6918 ( .C1(n12160), .C2(n2927), .B(n3017), .A(n11070), .ZN(n11067)
         );
  aoi21d1 U6919 ( .B1(images_bus[442]), .B2(n6557), .A(n11071), .ZN(n11065) );
  oai311d1 U6920 ( .C1(n9500), .C2(n11072), .C3(n11073), .A(n11074), .B(n11075), .ZN(n11063) );
  oai21d1 U6921 ( .B1(n10373), .B2(n9500), .A(n11076), .ZN(n11075) );
  aoi21d1 U6922 ( .B1(n3010), .B2(n2938), .A(n7194), .ZN(n10373) );
  oai321d1 U6925 ( .C1(n4795), .C2(n11080), .C3(n9512), .B1(n8746), .B2(n11081), .A(n11082), .ZN(n11079) );
  aoi21d1 U6928 ( .B1(n6598), .B2(n9504), .A(n4791), .ZN(n8746) );
  aoi321d1 U6930 ( .C1(n11083), .C2(n10370), .C3(images_bus[454]), .B1(n10235), 
        .B2(n11084), .A(n11085), .ZN(n11080) );
  oai31d1 U6931 ( .B1(n11086), .B2(n7313), .B3(n8756), .A(n9511), .ZN(n11085)
         );
  aon211d1 U6933 ( .C1(n7316), .C2(n6818), .B(n7315), .A(n11088), .ZN(n11086)
         );
  oai211d1 U6934 ( .C1(n11089), .C2(n2999), .A(n11090), .B(n11091), .ZN(n11084) );
  oai211d1 U6935 ( .C1(n10247), .C2(n7319), .A(n11092), .B(n3003), .ZN(n11091)
         );
  oaim21d1 U6937 ( .B1(n11088), .B2(n6818), .A(images_bus[459]), .ZN(n11092)
         );
  oai322d1 U6940 ( .C1(n9597), .C2(n11096), .C3(n10366), .A1(n10366), .A2(
        n11097), .B1(n2958), .B2(n11099), .ZN(n11095) );
  aon211d1 U6942 ( .C1(images_bus[466]), .C2(n10258), .B(n9597), .A(n11100), 
        .ZN(n11097) );
  aoi321d1 U6943 ( .C1(n2974), .C2(n11101), .C3(n7326), .B1(n2988), .B2(n11103), .A(n11104), .ZN(n11096) );
  oan211d1 U6944 ( .C1(n9526), .C2(n11105), .B(n11106), .A(n2986), .ZN(n11104)
         );
  aon211d1 U6946 ( .C1(n6212), .C2(n7333), .B(n10361), .A(n11108), .ZN(n11105)
         );
  oai321d1 U6950 ( .C1(n11109), .C2(n9543), .C3(n10271), .B1(n9538), .B2(
        n11110), .A(n11111), .ZN(n11101) );
  aoi22d1 U6951 ( .A1(n2975), .A2(n11113), .B1(n9533), .B2(n11114), .ZN(n11111) );
  oai21d1 U6952 ( .B1(n2984), .B2(n6982), .A(n2983), .ZN(n9533) );
  oai21d1 U6953 ( .B1(n11115), .B2(n10357), .A(n11116), .ZN(n11113) );
  oai211d1 U6954 ( .C1(n6425), .C2(n10357), .A(n9543), .B(n11117), .ZN(n11116)
         );
  aoi31d1 U6956 ( .B1(n11120), .B2(n2846), .B3(n2842), .A(n11122), .ZN(n11119)
         );
  aoi21d1 U6959 ( .B1(n7335), .B2(images_bus[480]), .A(n8796), .ZN(n8832) );
  oai22d1 U6960 ( .A1(n2913), .A2(n11124), .B1(n11125), .B2(n7337), .ZN(n11118) );
  aoi321d1 U6961 ( .C1(n2858), .C2(n5221), .C3(n11126), .B1(n9591), .B2(n11127), .A(n11128), .ZN(n11125) );
  aoi211d1 U6962 ( .C1(n11129), .C2(n11126), .A(n12125), .B(n11124), .ZN(
        n11128) );
  oai322d1 U6963 ( .C1(n11130), .C2(n11131), .C3(n11132), .A1(n11133), .A2(
        n2863), .B1(n2864), .B2(n11131), .ZN(n11127) );
  aoi322d1 U6964 ( .C1(n9584), .C2(n5968), .C3(n2862), .A1(n8005), .A2(n11134), 
        .B1(n11135), .B2(n2860), .ZN(n11133) );
  oan211d1 U6966 ( .C1(n2871), .C2(n6817), .B(n11137), .A(n11138), .ZN(n11135)
         );
  oai22d1 U6967 ( .A1(n11139), .A2(n11140), .B1(n2816), .B2(n10352), .ZN(
        n11134) );
  aoi21d1 U6968 ( .B1(n11142), .B2(images_bus[492]), .A(n8828), .ZN(n10352) );
  aoi321d1 U6969 ( .C1(n9562), .C2(n11143), .C3(images_bus[492]), .B1(n8006), 
        .B2(n11144), .A(n11145), .ZN(n11139) );
  oai21d1 U6970 ( .B1(n9562), .B2(n11146), .A(n11147), .ZN(n11145) );
  aon211d1 U6973 ( .C1(images_bus[494]), .C2(n8810), .B(n2881), .A(n11150), 
        .ZN(n11146) );
  oai322d1 U6975 ( .C1(n7050), .C2(n11151), .C3(n2885), .A1(n11153), .A2(
        n10349), .B1(n10322), .B2(n11154), .ZN(n11144) );
  aon211d1 U6976 ( .C1(images_bus[498]), .C2(n11155), .B(n11156), .A(n11157), 
        .ZN(n11154) );
  oai21d1 U6977 ( .B1(n11151), .B2(n7050), .A(images_bus[497]), .ZN(n11157) );
  or02d0 U6978 ( .A1(n4920), .A2(n11155), .Z(n10349) );
  aoi221d1 U6979 ( .B1(n11158), .B2(n11159), .C1(n11160), .C2(n2908), .A(
        n11162), .ZN(n11153) );
  oan211d1 U6980 ( .C1(n11163), .C2(n2891), .B(n11164), .A(n10348), .ZN(n11162) );
  aon211d1 U6982 ( .C1(images_bus[502]), .C2(n9578), .B(n2891), .A(n11167), 
        .ZN(n11164) );
  aoi322d1 U6983 ( .C1(n9581), .C2(n11168), .C3(n2889), .A1(n2887), .A2(n11170), .B1(n9577), .B2(n11171), .ZN(n11163) );
  oai22d1 U6984 ( .A1(n2896), .A2(n11172), .B1(n2902), .B2(n11174), .ZN(n11171) );
  oai31d1 U6986 ( .B1(n10343), .B2(n10346), .B3(n11176), .A(n11177), .ZN(
        n11170) );
  aoi31d1 U6987 ( .B1(n2900), .B2(N15618), .B3(n11178), .A(n11179), .ZN(n11177) );
  oan211d1 U6989 ( .C1(n11176), .C2(n12152), .B(images_bus[509]), .A(n10341), 
        .ZN(n11178) );
  or02d0 U6991 ( .A1(n11172), .A2(n6654), .Z(n11174) );
  aoi21d1 U6992 ( .B1(n11168), .B2(images_bus[504]), .A(n5320), .ZN(n11172) );
  aoim21d1 U6993 ( .B1(n12152), .B2(n11181), .A(n11182), .ZN(n10346) );
  oaim21d1 U6997 ( .B1(n11167), .B2(images_bus[502]), .A(images_bus[503]), 
        .ZN(n11168) );
  oai21d1 U6998 ( .B1(n2814), .B2(n6508), .A(n4297), .ZN(n11167) );
  aon211d1 U7000 ( .C1(N15554), .C2(n10329), .B(n6979), .A(n2894), .ZN(n10333)
         );
  oan211d1 U7001 ( .C1(n2904), .C2(n6508), .B(N15474), .A(n2814), .ZN(n11160)
         );
  aon211d1 U7003 ( .C1(images_bus[497]), .C2(n11185), .B(n6723), .A(
        images_bus[499]), .ZN(n11158) );
  aoi21d1 U7007 ( .B1(n11150), .B2(images_bus[494]), .A(n5894), .ZN(n11151) );
  oai21d1 U7008 ( .B1(n2816), .B2(n6553), .A(images_bus[493]), .ZN(n11150) );
  oai21d1 U7015 ( .B1(n11138), .B2(n6817), .A(images_bus[491]), .ZN(n11143) );
  oan211d1 U7016 ( .C1(n5968), .C2(n11188), .B(images_bus[488]), .A(n12166), 
        .ZN(n11138) );
  oan211d1 U7021 ( .C1(n10296), .C2(n9584), .B(images_bus[486]), .A(n9590), 
        .ZN(n11132) );
  oai21d1 U7022 ( .B1(n11190), .B2(n7115), .A(n11191), .ZN(n9584) );
  oan211d1 U7024 ( .C1(n5221), .C2(n11192), .B(images_bus[484]), .A(n4633), 
        .ZN(n11131) );
  aoi21d1 U7028 ( .B1(n11194), .B2(images_bus[484]), .A(n9594), .ZN(n11129) );
  aoi21d1 U7030 ( .B1(n11120), .B2(images_bus[480]), .A(n5715), .ZN(n11124) );
  oai21d1 U7031 ( .B1(n12161), .B2(n11123), .A(images_bus[479]), .ZN(n11120)
         );
  aon211d1 U7035 ( .C1(images_bus[474]), .C2(n8781), .B(n8774), .A(n11195), 
        .ZN(n11110) );
  oai21d1 U7038 ( .B1(n2977), .B2(n8774), .A(n2976), .ZN(n9536) );
  aon211d1 U7043 ( .C1(n10280), .C2(n6155), .B(n9542), .A(n2813), .ZN(n11109)
         );
  aoi21d1 U7045 ( .B1(n11117), .B2(n6425), .A(n2819), .ZN(n11123) );
  oaim21d1 U7046 ( .B1(n11195), .B2(images_bus[474]), .A(images_bus[475]), 
        .ZN(n11117) );
  oaim21d1 U7047 ( .B1(n11114), .B2(images_bus[472]), .A(images_bus[473]), 
        .ZN(n11195) );
  oaim21d1 U7048 ( .B1(n11108), .B2(n6212), .A(images_bus[471]), .ZN(n11114)
         );
  oaim21d1 U7049 ( .B1(n11103), .B2(n6512), .A(images_bus[469]), .ZN(n11108)
         );
  oaim21d1 U7050 ( .B1(n11100), .B2(images_bus[466]), .A(images_bus[467]), 
        .ZN(n11103) );
  aoi31d1 U7054 ( .B1(n11200), .B2(n10367), .B3(n2994), .A(n11201), .ZN(n11089) );
  oan211d1 U7055 ( .C1(n12156), .C2(n2995), .B(n2998), .A(n11203), .ZN(n11201)
         );
  oai211d1 U7056 ( .C1(n2967), .C2(n7057), .A(n2993), .B(n2992), .ZN(n10367)
         );
  oai21d1 U7058 ( .B1(n12156), .B2(n11203), .A(images_bus[463]), .ZN(n11200)
         );
  aoim21d1 U7059 ( .B1(n11204), .B2(n6555), .A(n4397), .ZN(n11203) );
  aoi21d1 U7062 ( .B1(n11088), .B2(n6818), .A(n5126), .ZN(n11204) );
  aon211d1 U7064 ( .C1(images_bus[455]), .C2(n11205), .B(n7117), .A(
        images_bus[457]), .ZN(n11088) );
  oai21d1 U7068 ( .B1(n3004), .B2(n7117), .A(n2950), .ZN(n11087) );
  oai21d1 U7069 ( .B1(n12141), .B2(n11081), .A(images_bus[453]), .ZN(n11083)
         );
  aoim21d1 U7070 ( .B1(n11072), .B2(n6894), .A(n5231), .ZN(n11081) );
  aoi31d1 U7072 ( .B1(n3010), .B2(n11206), .B3(n2938), .A(n11207), .ZN(n11073)
         );
  oai211d1 U7075 ( .C1(n3008), .C2(n6894), .A(n3009), .B(n2939), .ZN(n11206)
         );
  aoi21d1 U7077 ( .B1(n11076), .B2(images_bus[448]), .A(n5727), .ZN(n11072) );
  oai21d1 U7078 ( .B1(n11070), .B2(n12160), .A(images_bus[447]), .ZN(n11076)
         );
  aoi21d1 U7079 ( .B1(n11061), .B2(images_bus[444]), .A(n2915), .ZN(n11070) );
  aon211d1 U7081 ( .C1(n11058), .C2(n5354), .B(n6658), .A(images_bus[443]), 
        .ZN(n11061) );
  aon211d1 U7085 ( .C1(images_bus[437]), .C2(n11211), .B(n6218), .A(
        images_bus[439]), .ZN(n11055) );
  oai21d1 U7089 ( .B1(n3111), .B2(n6218), .A(n3094), .ZN(n11049) );
  aoi21d1 U7091 ( .B1(images_bus[431]), .B2(n11213), .A(n8712), .ZN(n11042) );
  aoi21d1 U7092 ( .B1(n7062), .B2(n11047), .A(n5600), .ZN(n8712) );
  oan211d1 U7093 ( .C1(n3093), .C2(n6519), .B(n3114), .A(n11212), .ZN(n11041)
         );
  aoi21d1 U7094 ( .B1(n11048), .B2(images_bus[434]), .A(n5003), .ZN(n11212) );
  aon211d1 U7095 ( .C1(images_bus[431]), .C2(n11213), .B(n12119), .A(
        images_bus[433]), .ZN(n11048) );
  aon211d1 U7097 ( .C1(images_bus[427]), .C2(n11032), .B(n12142), .A(
        images_bus[429]), .ZN(n11040) );
  or02d0 U7098 ( .A1(n11027), .A2(n6826), .Z(n11032) );
  oan211d1 U7103 ( .C1(n5980), .C2(n11021), .B(images_bus[424]), .A(n5617), 
        .ZN(n11027) );
  oai21d1 U7106 ( .B1(n11017), .B2(n12140), .A(images_bus[421]), .ZN(n11023)
         );
  aoi21d1 U7107 ( .B1(n11018), .B2(images_bus[418]), .A(n5235), .ZN(n11017) );
  oaim21d1 U7108 ( .B1(n11011), .B2(images_bus[416]), .A(images_bus[417]), 
        .ZN(n11018) );
  aoim21d1 U7109 ( .B1(n7939), .B2(n7121), .A(n9468), .ZN(n9464) );
  oai21d1 U7112 ( .B1(n11215), .B2(n6160), .A(images_bus[415]), .ZN(n11011) );
  oai21d1 U7113 ( .B1(n3043), .B2(n7205), .A(n3038), .ZN(n8682) );
  oan211d1 U7115 ( .C1(n3128), .C2(n6160), .B(n3031), .A(n11215), .ZN(n11005)
         );
  aoi21d1 U7116 ( .B1(n11004), .B2(n6437), .A(n3129), .ZN(n11215) );
  oai21d1 U7119 ( .B1(n12150), .B2(n9453), .A(n3227), .ZN(n10388) );
  oaim21d1 U7120 ( .B1(n6659), .B2(n11217), .A(images_bus[411]), .ZN(n11004)
         );
  aon211d1 U7121 ( .C1(n6424), .C2(n6659), .B(n8658), .A(n11217), .ZN(n11001)
         );
  oai21d1 U7122 ( .B1(n10998), .B2(n6993), .A(images_bus[409]), .ZN(n11217) );
  aoim21d1 U7125 ( .B1(n6406), .B2(n6581), .A(n11218), .ZN(n10999) );
  aoi21d1 U7128 ( .B1(n5552), .B2(images_bus[408]), .A(n6421), .ZN(n6581) );
  aoim21d1 U7129 ( .B1(n10997), .B2(n6225), .A(n5806), .ZN(n10998) );
  oan211d1 U7131 ( .C1(n5034), .C2(n10991), .B(images_bus[404]), .A(n4302), 
        .ZN(n10997) );
  oai21d1 U7132 ( .B1(images_bus[404]), .B2(n9438), .A(n6407), .ZN(n8837) );
  oan211d1 U7139 ( .C1(n5906), .C2(n11221), .B(images_bus[400]), .A(n5506), 
        .ZN(n10988) );
  aoi21d1 U7143 ( .B1(n10980), .B2(images_bus[396]), .A(n12171), .ZN(n10983)
         );
  oai21d1 U7145 ( .B1(n3195), .B2(n7066), .A(n3199), .ZN(n7235) );
  oai21d1 U7148 ( .B1(n3191), .B2(n6558), .A(n3186), .ZN(n10138) );
  oaim21d1 U7149 ( .B1(n10977), .B2(images_bus[394]), .A(images_bus[395]), 
        .ZN(n10980) );
  oai21d1 U7152 ( .B1(n10975), .B2(n7127), .A(images_bus[393]), .ZN(n10977) );
  oan211d1 U7154 ( .C1(n4649), .C2(n11223), .B(images_bus[390]), .A(n5982), 
        .ZN(n10975) );
  aon211d1 U7160 ( .C1(images_bus[385]), .C2(n10965), .B(n12124), .A(
        images_bus[387]), .ZN(n10967) );
  oai21d1 U7162 ( .B1(n10955), .B2(n6162), .A(images_bus[383]), .ZN(n10961) );
  aoi21d1 U7163 ( .B1(n10946), .B2(images_bus[380]), .A(n3138), .ZN(n10955) );
  oaim21d1 U7165 ( .B1(n10940), .B2(n6664), .A(images_bus[379]), .ZN(n10946)
         );
  oai21d1 U7166 ( .B1(n10950), .B2(n6997), .A(images_bus[377]), .ZN(n10940) );
  aoi21d1 U7168 ( .B1(n10944), .B2(images_bus[374]), .A(n5818), .ZN(n10950) );
  aon211d1 U7169 ( .C1(images_bus[371]), .C2(n11224), .B(n6525), .A(
        images_bus[373]), .ZN(n10944) );
  aoi21d1 U7172 ( .B1(images_bus[382]), .B2(n11225), .A(n7211), .ZN(n10954) );
  aon211d1 U7178 ( .C1(images_bus[367]), .C2(n11226), .B(n7067), .A(
        images_bus[369]), .ZN(n10936) );
  aoi21d1 U7184 ( .B1(n11230), .B2(images_bus[364]), .A(n4419), .ZN(n10934) );
  aon211d1 U7186 ( .C1(images_bus[364]), .C2(n11231), .B(n4601), .A(n11230), 
        .ZN(n10925) );
  oai21d1 U7187 ( .B1(n10923), .B2(n6838), .A(images_bus[363]), .ZN(n11230) );
  aoim21d1 U7188 ( .B1(n10919), .B2(n7133), .A(n12165), .ZN(n10923) );
  oan211d1 U7190 ( .C1(n4653), .C2(n11232), .B(images_bus[358]), .A(n5988), 
        .ZN(n10919) );
  aoi21d1 U7192 ( .B1(n3321), .B2(n6368), .A(n10915), .ZN(n10916) );
  aoi21d1 U7193 ( .B1(n6908), .B2(n10911), .A(n5249), .ZN(n10915) );
  oai21d1 U7195 ( .B1(n10907), .B2(n7222), .A(images_bus[353]), .ZN(n10911) );
  aoi21d1 U7196 ( .B1(n10906), .B2(images_bus[350]), .A(n6097), .ZN(n10907) );
  aon211d1 U7198 ( .C1(images_bus[347]), .C2(n11233), .B(n6445), .A(
        images_bus[349]), .ZN(n10906) );
  aon211d1 U7200 ( .C1(images_bus[346]), .C2(n10898), .B(n4915), .A(n8579), 
        .ZN(n10900) );
  aon211d1 U7202 ( .C1(images_bus[343]), .C2(n10897), .B(n6998), .A(
        images_bus[345]), .ZN(n10898) );
  aon211d1 U7204 ( .C1(images_bus[339]), .C2(n11234), .B(n6529), .A(
        images_bus[341]), .ZN(n10893) );
  aoi21d1 U7207 ( .B1(n3383), .B2(n6529), .A(n6251), .ZN(n10886) );
  oai21d1 U7209 ( .B1(n10881), .B2(n7069), .A(images_bus[337]), .ZN(n10879) );
  aoi21d1 U7210 ( .B1(n10884), .B2(images_bus[334]), .A(n5927), .ZN(n10881) );
  oai21d1 U7211 ( .B1(n10873), .B2(n6562), .A(images_bus[333]), .ZN(n10884) );
  oan211d1 U7212 ( .C1(n5633), .C2(n11235), .B(images_bus[330]), .A(n5156), 
        .ZN(n10873) );
  oan211d1 U7214 ( .C1(n4663), .C2(n11236), .B(images_bus[326]), .A(n6004), 
        .ZN(n10868) );
  oai21d1 U7217 ( .B1(n10859), .B2(n6919), .A(images_bus[323]), .ZN(n10864) );
  oan211d1 U7218 ( .C1(n6098), .C2(n11237), .B(images_bus[320]), .A(n5737), 
        .ZN(n10859) );
  oaim21d1 U7228 ( .B1(n11241), .B2(images_bus[316]), .A(images_bus[317]), 
        .ZN(n10851) );
  aon211d1 U7229 ( .C1(images_bus[316]), .C2(n5418), .B(n5420), .A(n11241), 
        .ZN(n10848) );
  oai21d1 U7230 ( .B1(n3485), .B2(n6675), .A(images_bus[315]), .ZN(n11241) );
  aon211d1 U7237 ( .C1(images_bus[311]), .C2(n10840), .B(n7006), .A(
        images_bus[313]), .ZN(n10843) );
  or02d0 U7239 ( .A1(n10835), .A2(n6240), .Z(n10840) );
  aoi21d1 U7240 ( .B1(n6531), .B2(n10834), .A(n4307), .ZN(n10835) );
  oai21d1 U7241 ( .B1(n10831), .B2(n6752), .A(images_bus[307]), .ZN(n10834) );
  aoim21d1 U7243 ( .B1(n10827), .B2(n7072), .A(n5531), .ZN(n10831) );
  oan211d1 U7245 ( .C1(n4436), .C2(n10830), .B(images_bus[302]), .A(n5931), 
        .ZN(n10827) );
  aoi21d1 U7248 ( .B1(n10824), .B2(images_bus[298]), .A(n5164), .ZN(n10819) );
  oaim21d1 U7249 ( .B1(n10816), .B2(images_bus[296]), .A(images_bus[297]), 
        .ZN(n10824) );
  oai21d1 U7252 ( .B1(n10814), .B2(n12153), .A(images_bus[295]), .ZN(n10816)
         );
  aoi21d1 U7253 ( .B1(n10811), .B2(images_bus[292]), .A(n4675), .ZN(n10814) );
  oai21d1 U7254 ( .B1(n10805), .B2(n12122), .A(images_bus[291]), .ZN(n10811)
         );
  aoim21d1 U7255 ( .B1(n10804), .B2(n7237), .A(n5738), .ZN(n10805) );
  aoi21d1 U7258 ( .B1(n10794), .B2(images_bus[286]), .A(n6100), .ZN(n10804) );
  oai21d1 U7259 ( .B1(n10801), .B2(n12149), .A(images_bus[285]), .ZN(n10794)
         );
  aon211d1 U7261 ( .C1(images_bus[280]), .C2(n10791), .B(n5410), .A(
        images_bus[282]), .ZN(n10790) );
  oai21d1 U7263 ( .B1(n10786), .B2(n6242), .A(images_bus[279]), .ZN(n10791) );
  aoi21d1 U7264 ( .B1(n10779), .B2(images_bus[276]), .A(n4311), .ZN(n10786) );
  oai21d1 U7265 ( .B1(n11243), .B2(n6753), .A(images_bus[275]), .ZN(n10779) );
  or02d0 U7272 ( .A1(n4465), .A2(n4456), .Z(n9254) );
  aon211d1 U7273 ( .C1(n11245), .C2(n7762), .B(n11246), .A(n9250), .ZN(n10771)
         );
  aoi21d1 U7276 ( .B1(n11245), .B2(images_bus[272]), .A(n5540), .ZN(n11243) );
  aon211d1 U7278 ( .C1(images_bus[269]), .C2(n11247), .B(n6305), .A(
        images_bus[271]), .ZN(n11245) );
  aoi31d1 U7280 ( .B1(n10774), .B2(n7760), .B3(images_bus[268]), .A(n8484), 
        .ZN(n10770) );
  aon211d1 U7281 ( .C1(images_bus[265]), .C2(n10768), .B(n6849), .A(
        images_bus[267]), .ZN(n10774) );
  oai21d1 U7286 ( .B1(n10759), .B2(n6388), .A(images_bus[263]), .ZN(n10765) );
  aoi21d1 U7287 ( .B1(n10763), .B2(images_bus[260]), .A(n4689), .ZN(n10759) );
  oaim21d1 U7288 ( .B1(n10761), .B2(images_bus[258]), .A(images_bus[259]), 
        .ZN(n10763) );
  aon211d1 U7293 ( .C1(images_bus[255]), .C2(n10752), .B(n7240), .A(
        images_bus[257]), .ZN(n10761) );
  oai21d1 U7296 ( .B1(n10750), .B2(n6469), .A(images_bus[253]), .ZN(n10748) );
  aoi21d1 U7298 ( .B1(n10742), .B2(images_bus[250]), .A(n4948), .ZN(n10750) );
  oaim21d1 U7303 ( .B1(n10740), .B2(images_bus[248]), .A(images_bus[249]), 
        .ZN(n10742) );
  aon211d1 U7304 ( .C1(images_bus[245]), .C2(n11254), .B(n6246), .A(
        images_bus[247]), .ZN(n10740) );
  oan211d1 U7310 ( .C1(n5542), .C2(n10731), .B(images_bus[242]), .A(n5063), 
        .ZN(n10738) );
  oaim21d1 U7313 ( .B1(n10723), .B2(images_bus[238]), .A(images_bus[239]), 
        .ZN(n10724) );
  aon211d1 U7314 ( .C1(images_bus[235]), .C2(n10720), .B(n6567), .A(
        images_bus[237]), .ZN(n10723) );
  oai21d1 U7317 ( .B1(n10713), .B2(n12118), .A(images_bus[233]), .ZN(n10718)
         );
  aoim21d1 U7320 ( .B1(n10715), .B2(n6389), .A(n6025), .ZN(n10713) );
  oan211d1 U7323 ( .C1(n5268), .C2(n11255), .B(n6621), .A(n4691), .ZN(n10715)
         );
  oai21d1 U7330 ( .B1(n10710), .B2(n7242), .A(images_bus[225]), .ZN(n10711) );
  aoi21d1 U7331 ( .B1(n10704), .B2(images_bus[222]), .A(n6115), .ZN(n10710) );
  oai21d1 U7333 ( .B1(n10702), .B2(n6475), .A(images_bus[221]), .ZN(n10704) );
  oan211d1 U7335 ( .C1(n5431), .C2(n11256), .B(n6682), .A(n4951), .ZN(n10702)
         );
  aoi21d1 U7339 ( .B1(n10696), .B2(images_bus[214]), .A(n5839), .ZN(n10697) );
  oaim21d1 U7340 ( .B1(n10689), .B2(images_bus[212]), .A(images_bus[213]), 
        .ZN(n10696) );
  oaim21d1 U7341 ( .B1(n10690), .B2(images_bus[210]), .A(images_bus[211]), 
        .ZN(n10689) );
  oai21d1 U7342 ( .B1(n10687), .B2(n7079), .A(images_bus[209]), .ZN(n10690) );
  aoi21d1 U7344 ( .B1(n6324), .B2(n11258), .A(n5944), .ZN(n10687) );
  aoi31d1 U7349 ( .B1(n10683), .B2(n11258), .B3(n3878), .A(n5186), .ZN(n10679)
         );
  oai21d1 U7351 ( .B1(n11260), .B2(n6571), .A(images_bus[205]), .ZN(n11258) );
  aoi21d1 U7352 ( .B1(n10678), .B2(n6861), .A(n5186), .ZN(n11260) );
  oai21d1 U7353 ( .B1(n11261), .B2(n7155), .A(images_bus[201]), .ZN(n10678) );
  aoi21d1 U7354 ( .B1(images_bus[198]), .B2(n10673), .A(n6038), .ZN(n11261) );
  aon211d1 U7355 ( .C1(images_bus[195]), .C2(n11262), .B(n6628), .A(n4698), 
        .ZN(n10673) );
  aon211d1 U7357 ( .C1(images_bus[191]), .C2(n11263), .B(n7243), .A(
        images_bus[193]), .ZN(n10671) );
  oai21d1 U7359 ( .B1(n3906), .B2(n6481), .A(images_bus[189]), .ZN(n10667) );
  aon211d1 U7361 ( .C1(images_bus[185]), .C2(n10653), .B(n6683), .A(n4958), 
        .ZN(n11264) );
  oaim21d1 U7364 ( .B1(n10651), .B2(images_bus[182]), .A(images_bus[183]), 
        .ZN(n10650) );
  aon211d1 U7365 ( .C1(images_bus[179]), .C2(n11265), .B(n12145), .A(
        images_bus[181]), .ZN(n10651) );
  aon211d1 U7368 ( .C1(images_bus[175]), .C2(n11267), .B(n7081), .A(
        images_bus[177]), .ZN(n11266) );
  oai21d1 U7371 ( .B1(n10642), .B2(n6572), .A(images_bus[173]), .ZN(n11268) );
  aoim21d1 U7373 ( .B1(n10635), .B2(n6866), .A(n5189), .ZN(n10642) );
  aoi21d1 U7375 ( .B1(n10633), .B2(images_bus[168]), .A(n5676), .ZN(n10635) );
  oai21d1 U7378 ( .B1(n10629), .B2(n6395), .A(images_bus[167]), .ZN(n10633) );
  aoi21d1 U7380 ( .B1(n10628), .B2(images_bus[164]), .A(n4703), .ZN(n10629) );
  aon211d1 U7381 ( .C1(images_bus[161]), .C2(n11269), .B(n6938), .A(
        images_bus[163]), .ZN(n10628) );
  aon211d1 U7383 ( .C1(images_bus[157]), .C2(n11270), .B(n6185), .A(
        images_bus[159]), .ZN(n10624) );
  oaim21d1 U7386 ( .B1(n10620), .B2(images_bus[154]), .A(images_bus[155]), 
        .ZN(n10619) );
  oai21d1 U7387 ( .B1(n10615), .B2(n7023), .A(images_bus[153]), .ZN(n10620) );
  aoi21d1 U7390 ( .B1(n10611), .B2(images_bus[150]), .A(n5851), .ZN(n10615) );
  aon211d1 U7392 ( .C1(images_bus[146]), .C2(n10607), .B(n5098), .A(n6544), 
        .ZN(n11272) );
  aon211d1 U7393 ( .C1(images_bus[143]), .C2(n3987), .B(n7093), .A(
        images_bus[145]), .ZN(n10607) );
  aon211d1 U7396 ( .C1(n5090), .C2(n4027), .B(n5952), .A(n4053), .ZN(n10604)
         );
  oai21d1 U7401 ( .B1(n11274), .B2(n5074), .A(images_bus[139]), .ZN(n10598) );
  oan211d1 U7402 ( .C1(n5194), .C2(n10599), .B(images_bus[140]), .A(n4491), 
        .ZN(n11274) );
  aoi21d1 U7404 ( .B1(n10595), .B2(images_bus[136]), .A(n5684), .ZN(n10596) );
  aon211d1 U7405 ( .C1(images_bus[133]), .C2(n11276), .B(n6397), .A(
        images_bus[135]), .ZN(n10595) );
  aoi21d1 U7408 ( .B1(n10590), .B2(images_bus[130]), .A(n5281), .ZN(n10592) );
  oai21d1 U7409 ( .B1(n10586), .B2(n7245), .A(images_bus[129]), .ZN(n10590) );
  aoi21d1 U7410 ( .B1(n10583), .B2(images_bus[126]), .A(n6133), .ZN(n10586) );
  oai21d1 U7412 ( .B1(n10580), .B2(n6488), .A(images_bus[125]), .ZN(n10583) );
  aoi21d1 U7415 ( .B1(n10579), .B2(images_bus[122]), .A(n4965), .ZN(n10580) );
  aon211d1 U7416 ( .C1(images_bus[119]), .C2(n11278), .B(n7034), .A(
        images_bus[121]), .ZN(n10579) );
  aon211d1 U7421 ( .C1(images_bus[115]), .C2(n11280), .B(n12143), .A(
        images_bus[117]), .ZN(n11279) );
  oaim21d1 U7423 ( .B1(n10572), .B2(images_bus[112]), .A(images_bus[113]), 
        .ZN(n10571) );
  oai21d1 U7424 ( .B1(n10566), .B2(n6344), .A(images_bus[111]), .ZN(n10572) );
  aoim21d1 U7426 ( .B1(n10562), .B2(n6576), .A(n4493), .ZN(n10566) );
  oan211d1 U7428 ( .C1(n5689), .C2(n10565), .B(images_bus[106]), .A(n5203), 
        .ZN(n10562) );
  aon211d1 U7430 ( .C1(images_bus[101]), .C2(n11281), .B(n6400), .A(
        images_bus[103]), .ZN(n10561) );
  or02d0 U7431 ( .A1(n10554), .A2(n6639), .Z(n11281) );
  aoi21d1 U7436 ( .B1(n10559), .B2(images_bus[98]), .A(n5284), .ZN(n10554) );
  oai21d1 U7437 ( .B1(n10557), .B2(n7251), .A(images_bus[97]), .ZN(n10559) );
  aoi21d1 U7438 ( .B1(n10553), .B2(images_bus[94]), .A(n6138), .ZN(n10557) );
  aon211d1 U7441 ( .C1(images_bus[91]), .C2(n11282), .B(n12148), .A(
        images_bus[93]), .ZN(n10553) );
  oai21d1 U7445 ( .B1(n10546), .B2(n7042), .A(images_bus[89]), .ZN(n10548) );
  aoim21d1 U7448 ( .B1(n10545), .B2(n6268), .A(n5858), .ZN(n10546) );
  aoim21d1 U7450 ( .B1(n10543), .B2(n6548), .A(n4326), .ZN(n10545) );
  oan211d1 U7452 ( .C1(n5581), .C2(n11284), .B(images_bus[82]), .A(n5106), 
        .ZN(n10543) );
  aon211d1 U7455 ( .C1(images_bus[77]), .C2(n11285), .B(n6345), .A(
        images_bus[79]), .ZN(n10535) );
  oai21d1 U7468 ( .B1(n10525), .B2(n6882), .A(images_bus[75]), .ZN(n10530) );
  aoim21d1 U7469 ( .B1(n10522), .B2(n7182), .A(n5691), .ZN(n10525) );
  aoi21d1 U7470 ( .B1(n10524), .B2(images_bus[70]), .A(n6061), .ZN(n10522) );
  aon211d1 U7472 ( .C1(images_bus[67]), .C2(n10521), .B(n6641), .A(
        images_bus[69]), .ZN(n10524) );
  aoi31d1 U7475 ( .B1(n4199), .B2(n11288), .B3(n4195), .A(n11290), .ZN(n10515)
         );
  oaim21d1 U7476 ( .B1(n11290), .B2(images_bus[64]), .A(images_bus[65]), .ZN(
        n11288) );
  oai21d1 U7477 ( .B1(n10514), .B2(n6200), .A(images_bus[63]), .ZN(n11290) );
  oan211d1 U7478 ( .C1(n4974), .C2(n11291), .B(images_bus[60]), .A(n4222), 
        .ZN(n10514) );
  aon211d1 U7482 ( .C1(images_bus[55]), .C2(n10507), .B(n7045), .A(
        images_bus[57]), .ZN(n10509) );
  oai21d1 U7484 ( .B1(n4294), .B2(n6550), .A(n4331), .ZN(n10503) );
  aon211d1 U7486 ( .C1(images_bus[49]), .C2(n11292), .B(n12130), .A(
        images_bus[51]), .ZN(n10504) );
  aon211d1 U7488 ( .C1(images_bus[45]), .C2(n11293), .B(n6348), .A(
        images_bus[47]), .ZN(n10498) );
  aoi21d1 U7495 ( .B1(n10488), .B2(images_bus[42]), .A(n5205), .ZN(n10492) );
  aon211d1 U7498 ( .C1(images_bus[38]), .C2(n10484), .B(n6070), .A(
        images_bus[40]), .ZN(n11294) );
  oai21d1 U7499 ( .B1(n11295), .B2(n6646), .A(images_bus[37]), .ZN(n10484) );
  aoim21d1 U7500 ( .B1(n10477), .B2(n12120), .A(n5312), .ZN(n11295) );
  oan211d1 U7501 ( .C1(n6146), .C2(n10476), .B(images_bus[32]), .A(n5782), 
        .ZN(n10477) );
  aon211d1 U7507 ( .C1(images_bus[27]), .C2(n10467), .B(n6507), .A(
        images_bus[29]), .ZN(n10469) );
  oai21d1 U7509 ( .B1(n10462), .B2(n7047), .A(images_bus[25]), .ZN(n10464) );
  aon211d1 U7511 ( .C1(images_bus[20]), .C2(n10455), .B(n4342), .A(
        images_bus[22]), .ZN(n11296) );
  aon211d1 U7516 ( .C1(images_bus[17]), .C2(n10449), .B(n6813), .A(
        images_bus[19]), .ZN(n10455) );
  oai21d1 U7519 ( .B1(n11298), .B2(n6355), .A(images_bus[15]), .ZN(n10447) );
  aoi21d1 U7520 ( .B1(images_bus[12]), .B2(n4881), .A(n4608), .ZN(n11298) );
  aoi21d1 U7522 ( .B1(n6890), .B2(n10440), .A(n5220), .ZN(n10444) );
  aon211d1 U7525 ( .C1(images_bus[6]), .C2(n10437), .B(n6072), .A(
        images_bus[8]), .ZN(n11299) );
  oai21d1 U7526 ( .B1(n10435), .B2(n6653), .A(images_bus[5]), .ZN(n10437) );
  aoi21d1 U7527 ( .B1(n5785), .B2(images_bus[2]), .A(n5315), .ZN(n10435) );
  aor31d1 U7533 ( .B1(N8001), .B2(n11302), .B3(N7997), .A(n2772), .Z(N26357)
         );
  oai211d1 U7535 ( .C1(n9645), .C2(n7574), .A(n11303), .B(images_bus[1]), .ZN(
        n11302) );
  aon211d1 U7537 ( .C1(n11306), .C2(images_bus[4]), .B(n9652), .A(n11304), 
        .ZN(n11305) );
  aoi22d1 U7539 ( .A1(n4854), .A2(n11307), .B1(n8894), .B2(n4871), .ZN(n11306)
         );
  oai211d1 U7540 ( .C1(n11308), .C2(n10441), .A(n9656), .B(n11309), .ZN(n11307) );
  aoi21d1 U7541 ( .B1(n4767), .B2(n11311), .A(n9657), .ZN(n11309) );
  oan211d1 U7549 ( .C1(n11314), .C2(n11315), .B(n4789), .A(n12164), .ZN(n11308) );
  oan211d1 U7552 ( .C1(n11316), .C2(n7588), .B(n4827), .A(n9661), .ZN(n11314)
         );
  aoi321d1 U7555 ( .C1(n4628), .C2(n11319), .C3(n9659), .B1(n4816), .B2(n4608), 
        .A(n10445), .ZN(n11316) );
  aon211d1 U7559 ( .C1(n11320), .C2(n11321), .B(n10453), .A(n9663), .ZN(n11319) );
  aoi21d1 U7560 ( .B1(n5964), .B2(n4604), .A(n6355), .ZN(n9663) );
  aoi211d1 U7565 ( .C1(n7468), .C2(n4575), .A(n4580), .B(n7471), .ZN(n11321)
         );
  aoi211d1 U7573 ( .C1(n7472), .C2(n11325), .A(n10452), .B(n11326), .ZN(n11320) );
  aoi31d1 U7574 ( .B1(n4392), .B2(n11327), .B3(n7478), .A(n4551), .ZN(n11326)
         );
  aoi22d1 U7586 ( .A1(n6273), .A2(n4365), .B1(n11330), .B2(n4357), .ZN(n7478)
         );
  oai211d1 U7589 ( .C1(n4369), .C2(n11330), .A(n11331), .B(n11297), .ZN(n11327) );
  aon211d1 U7594 ( .C1(n7484), .C2(n9684), .B(n11332), .A(n11333), .ZN(n11331)
         );
  oan211d1 U7598 ( .C1(n11337), .C2(n9696), .B(n11338), .A(n4280), .ZN(n11335)
         );
  oai21d1 U7607 ( .B1(n11342), .B2(n10478), .A(images_bus[32]), .ZN(n6668) );
  oai22d1 U7608 ( .A1(images_bus[33]), .A2(n6686), .B1(n11343), .B2(n4231), 
        .ZN(n11340) );
  aoim2m11d1 U7612 ( .C1(n8937), .C2(n11344), .B(n6687), .A(n11345), .ZN(
        n11343) );
  aon211d1 U7613 ( .C1(n11346), .C2(n11347), .B(n4238), .A(n6967), .ZN(n11345)
         );
  oai21d1 U7617 ( .B1(n11349), .B2(n11350), .A(n4275), .ZN(n11347) );
  oai21d1 U7618 ( .B1(n6702), .B2(n7458), .A(n9704), .ZN(n11350) );
  ora31d1 U7620 ( .B1(n11352), .B2(n6706), .B3(n11353), .A(n5788), .Z(n11349)
         );
  oai322d1 U7626 ( .C1(n6713), .C2(n11354), .C3(n5800), .A1(n6711), .A2(n11355), .B1(n6710), .B2(n11356), .ZN(n11353) );
  ora211d1 U7628 ( .C1(n11359), .C2(n9714), .A(n6714), .B(n11356), .Z(n11354)
         );
  aoi21d1 U7629 ( .B1(n5959), .B2(n4271), .A(n8204), .ZN(n6714) );
  nd13d1 U7632 ( .A1(n8204), .A2(n8197), .A3(N8536), .ZN(n8957) );
  oai21d1 U7637 ( .B1(n4229), .B2(n4255), .A(images_bus[47]), .ZN(n11361) );
  oai211d1 U7638 ( .C1(n11364), .C2(n4256), .A(n7517), .B(n11365), .ZN(n11360)
         );
  aoi22d1 U7639 ( .A1(n7454), .A2(n11366), .B1(n6721), .B2(n11367), .ZN(n11365) );
  oai21d1 U7644 ( .B1(n5110), .B2(n11369), .A(n7511), .ZN(n7517) );
  oai22d1 U7645 ( .A1(n8214), .A2(n8965), .B1(n11370), .B2(n10508), .ZN(n11369) );
  aoi211d1 U7667 ( .C1(n4261), .C2(n11376), .A(n11366), .B(n6725), .ZN(n11364)
         );
  aoim21d1 U7669 ( .B1(n11377), .B2(n8971), .A(n7045), .ZN(n8221) );
  aoi21d1 U7671 ( .B1(n4268), .B2(n11378), .A(n5459), .ZN(n11377) );
  aoi221d1 U7674 ( .B1(n4264), .B2(n11383), .C1(n6734), .C2(n11384), .A(n4265), 
        .ZN(n11382) );
  oai211d1 U7679 ( .C1(n8884), .C2(n8992), .A(n8115), .B(images_bus[61]), .ZN(
        n11383) );
  oai31d1 U7681 ( .B1(n11384), .B2(n7452), .B3(n11386), .A(n4146), .ZN(n11380)
         );
  aor221d1 U7694 ( .B1(n4188), .B2(n5298), .C1(n4191), .C2(n11388), .A(n11389), 
        .Z(n11386) );
  oan211d1 U7695 ( .C1(images_bus[65]), .C2(n11390), .B(images_bus[64]), .A(
        n5793), .ZN(n11389) );
  oai211d1 U7696 ( .C1(n11391), .C2(n5018), .A(images_bus[65]), .B(
        images_bus[66]), .ZN(n11388) );
  aoi31d1 U7700 ( .B1(n11392), .B2(n11393), .B3(n10423), .A(n11394), .ZN(
        n11391) );
  oai211d1 U7702 ( .C1(n11395), .C2(n9004), .A(images_bus[69]), .B(n11396), 
        .ZN(n11393) );
  oan211d1 U7703 ( .C1(n4148), .C2(n5815), .B(n9008), .A(n11398), .ZN(n11396)
         );
  aoi211d1 U7704 ( .C1(n4145), .C2(n11400), .A(n10527), .B(n5691), .ZN(n11398)
         );
  oai31d1 U7708 ( .B1(n11401), .B2(n6882), .B3(n11402), .A(n4152), .ZN(n11400)
         );
  aon211d1 U7712 ( .C1(n11403), .C2(n11404), .B(n7541), .A(n8249), .ZN(n11401)
         );
  oan211d1 U7718 ( .C1(n11406), .C2(n11407), .B(n5042), .A(n8251), .ZN(n11403)
         );
  aoi31d1 U7723 ( .B1(n11404), .B2(n5840), .B3(n11408), .A(n11409), .ZN(n11406) );
  aoi22d1 U7724 ( .A1(n6762), .A2(n11410), .B1(n7548), .B2(n11411), .ZN(n11408) );
  oai211d1 U7725 ( .C1(n11412), .C2(n6765), .A(images_bus[81]), .B(n4143), 
        .ZN(n11410) );
  oan211d1 U7728 ( .C1(n11414), .C2(n11415), .B(n4173), .A(n7551), .ZN(n11412)
         );
  oai21d1 U7729 ( .B1(n11416), .B2(n10544), .A(images_bus[82]), .ZN(n7551) );
  aoim31d1 U7735 ( .B1(n11287), .B2(images_bus[85]), .B3(n6768), .A(n11418), 
        .ZN(n7554) );
  oan211d1 U7736 ( .C1(images_bus[87]), .C2(n5859), .B(n6661), .A(n4161), .ZN(
        n11418) );
  oai22d1 U7737 ( .A1(n11419), .A2(n11287), .B1(n4161), .B2(n11420), .ZN(
        n11414) );
  aon211d1 U7738 ( .C1(n4169), .C2(n11421), .B(n11422), .A(n4171), .ZN(n11420)
         );
  aon211d1 U7743 ( .C1(n7564), .C2(n11424), .B(n8110), .A(n11425), .ZN(n11421)
         );
  aon211d1 U7749 ( .C1(n8105), .C2(n11426), .B(n11427), .A(n8104), .ZN(n11424)
         );
  oai211d1 U7750 ( .C1(n11428), .C2(n5874), .A(n5875), .B(n4144), .ZN(n11426)
         );
  aoi21d1 U7752 ( .B1(n5879), .B2(n4118), .A(n4119), .ZN(n5875) );
  aoim211d1 U7757 ( .C1(n5881), .C2(n11431), .A(n5878), .B(n11432), .ZN(n11428) );
  oan211d1 U7758 ( .C1(n11433), .C2(n11434), .B(n11435), .A(n5882), .ZN(n11432) );
  aoi311d1 U7763 ( .C1(n5886), .C2(n5895), .C3(n11436), .A(n11437), .B(n6783), 
        .ZN(n11433) );
  aon211d1 U7765 ( .C1(n5889), .C2(n11438), .B(n4114), .A(n11435), .ZN(n11437)
         );
  aoi21d1 U7769 ( .B1(n4745), .B2(n5895), .A(n11440), .ZN(n5889) );
  aoi21d1 U7770 ( .B1(images_bus[103]), .B2(n11441), .A(n4067), .ZN(n11436) );
  aon211d1 U7775 ( .C1(n4071), .C2(n11444), .B(n11439), .A(n8282), .ZN(n11441)
         );
  oai211d1 U7776 ( .C1(n11445), .C2(n6797), .A(n6656), .B(n4138), .ZN(n11444)
         );
  oai21d1 U7777 ( .B1(n5909), .B2(n5689), .A(n4111), .ZN(n6797) );
  oan211d1 U7783 ( .C1(n2790), .C2(n8290), .B(n11450), .A(n6803), .ZN(n11447)
         );
  oaim211d1 U7787 ( .C1(n4078), .C2(n11452), .A(n11450), .B(n6800), .ZN(n11451) );
  aoi22d1 U7788 ( .A1(n4493), .A2(n4079), .B1(n7442), .B2(n4078), .ZN(n6800)
         );
  oai222d1 U7790 ( .A1(n4083), .A2(n5026), .B1(n11453), .B2(n8297), .C1(n11454), .C2(n5923), .ZN(n11452) );
  aoi31d1 U7792 ( .B1(n4083), .B2(n11456), .B3(n4104), .A(n11457), .ZN(n11453)
         );
  oai211d1 U7793 ( .C1(n11458), .C2(n5017), .A(images_bus[113]), .B(n11454), 
        .ZN(n11456) );
  aoi211d1 U7795 ( .C1(n4085), .C2(n11459), .A(n5926), .B(n4084), .ZN(n11458)
         );
  aon211d1 U7800 ( .C1(n4099), .C2(n11461), .B(n11462), .A(n6821), .ZN(n11460)
         );
  oai21d1 U7805 ( .B1(n11463), .B2(n5030), .A(n7439), .ZN(n11461) );
  oai211d1 U7811 ( .C1(n7600), .C2(n6830), .A(n11465), .B(images_bus[119]), 
        .ZN(n11464) );
  aon211d1 U7812 ( .C1(n4094), .C2(n11467), .B(n11468), .A(n5024), .ZN(n11465)
         );
  aon211d1 U7814 ( .C1(n4966), .C2(n11469), .B(n6835), .A(n6831), .ZN(n11467)
         );
  aoi31d1 U7815 ( .B1(n4098), .B2(n3986), .B3(n4097), .A(n4965), .ZN(n6831) );
  oai311d1 U7820 ( .C1(n11471), .C2(n6649), .C3(n11468), .A(n3999), .B(n4098), 
        .ZN(n11469) );
  aon211d1 U7825 ( .C1(images_bus[127]), .C2(n11472), .B(n10587), .A(n4966), 
        .ZN(n11471) );
  aon211d1 U7827 ( .C1(n11473), .C2(n11474), .B(n3994), .A(n4001), .ZN(n11472)
         );
  aon211d1 U7831 ( .C1(n11477), .C2(images_bus[129]), .B(n5006), .A(n11478), 
        .ZN(n11474) );
  aoi22d1 U7833 ( .A1(n4004), .A2(n11479), .B1(n4006), .B2(n6946), .ZN(n11477)
         );
  oai211d1 U7834 ( .C1(n11480), .C2(n11277), .A(n11481), .B(n11482), .ZN(
        n11479) );
  aon211d1 U7835 ( .C1(n4014), .C2(n11483), .B(n11484), .A(n6648), .ZN(n11481)
         );
  oai211d1 U7838 ( .C1(n11485), .C2(n10593), .A(images_bus[133]), .B(n11480), 
        .ZN(n11483) );
  aoi211d1 U7840 ( .C1(n9098), .C2(n6051), .A(n6397), .B(n11486), .ZN(n11485)
         );
  aoi31d1 U7841 ( .B1(n11487), .B2(n8870), .B3(n11488), .A(n8320), .ZN(n11486)
         );
  aoi22d1 U7844 ( .A1(n4018), .A2(n11489), .B1(n4019), .B2(n5684), .ZN(n11488)
         );
  aon211d1 U7845 ( .C1(n11491), .C2(n11492), .B(n11493), .A(n11491), .ZN(
        n11489) );
  oai21d1 U7846 ( .B1(n5194), .B2(n11494), .A(n10603), .ZN(n11492) );
  oaim22d1 U7848 ( .A1(n11495), .A2(n5074), .B1(n11496), .B2(n4022), .ZN(
        n11494) );
  aoi211d1 U7854 ( .C1(n4025), .C2(n11497), .A(n11496), .B(n4491), .ZN(n11495)
         );
  oai211d1 U7855 ( .C1(n11498), .C2(n5076), .A(n11499), .B(n5077), .ZN(n11497)
         );
  oai21d1 U7856 ( .B1(n11500), .B2(n7626), .A(n4026), .ZN(n11499) );
  oai21d1 U7861 ( .B1(images_bus[145]), .B2(n10609), .A(images_bus[144]), .ZN(
        n7626) );
  aoi31d1 U7862 ( .B1(n11498), .B2(n5570), .B3(n11501), .A(n5084), .ZN(n11500)
         );
  nd13d1 U7863 ( .A1(n10609), .A2(N9921), .A3(n11502), .ZN(n5084) );
  aoi221d1 U7867 ( .B1(n5088), .B2(n11504), .C1(n4049), .C2(n11505), .A(n5090), 
        .ZN(n11501) );
  oaim211d1 U7869 ( .C1(n8096), .C2(n8095), .A(n3993), .B(n11507), .ZN(n11505)
         );
  aoi221d1 U7870 ( .B1(n4035), .B2(n11508), .C1(n7633), .C2(n11509), .A(n7635), 
        .ZN(n11507) );
  oai211d1 U7873 ( .C1(n11511), .C2(n10414), .A(n7639), .B(n5783), .ZN(n11509)
         );
  nd13d1 U7874 ( .A1(n8340), .A2(n4034), .A3(n10617), .ZN(n7639) );
  aoi211d1 U7878 ( .C1(n4042), .C2(n11513), .A(n11508), .B(n5103), .ZN(n11511)
         );
  oai21d1 U7879 ( .B1(images_bus[155]), .B2(n9847), .A(images_bus[153]), .ZN(
        n5103) );
  oai211d1 U7880 ( .C1(n11514), .C2(n8343), .A(n5442), .B(n3992), .ZN(n11513)
         );
  aoi211d1 U7887 ( .C1(n11516), .C2(n7647), .A(n5112), .B(n9122), .ZN(n11514)
         );
  aoi22d1 U7894 ( .A1(n11517), .A2(n11518), .B1(n11519), .B2(n7650), .ZN(
        n11516) );
  aon211d1 U7896 ( .C1(n5120), .C2(n11520), .B(n7244), .A(n3968), .ZN(n11518)
         );
  oai211d1 U7900 ( .C1(n11521), .C2(n5123), .A(n5763), .B(n11517), .ZN(n11520)
         );
  oan211d1 U7903 ( .C1(n11522), .C2(n11523), .B(n3914), .A(n11524), .ZN(n11521) );
  or02d0 U7906 ( .A1(n11524), .A2(n10632), .Z(n11523) );
  aon211d1 U7907 ( .C1(n11525), .C2(n5128), .B(n5131), .A(images_bus[163]), 
        .ZN(n11522) );
  aoi21d1 U7909 ( .B1(n4703), .B2(n3921), .A(n6630), .ZN(n5128) );
  oan211d1 U7912 ( .C1(n11527), .C2(n5139), .B(n3919), .A(n11529), .ZN(n11525)
         );
  oan211d1 U7913 ( .C1(images_bus[167]), .C2(n5135), .B(n4711), .A(n5137), 
        .ZN(n11529) );
  aoi211d1 U7924 ( .C1(n11530), .C2(n3925), .A(n5994), .B(n7166), .ZN(n11527)
         );
  oai22d1 U7926 ( .A1(images_bus[169]), .A2(n5144), .B1(n11532), .B2(n3926), 
        .ZN(n8358) );
  aoi22d1 U7927 ( .A1(n3929), .A2(n11533), .B1(n3928), .B2(n7430), .ZN(n11532)
         );
  aor31d1 U7928 ( .B1(n3933), .B2(n4464), .B3(n11534), .A(n5189), .Z(n11533)
         );
  aon211d1 U7934 ( .C1(n5163), .C2(n11538), .B(n5155), .A(n5157), .ZN(n11537)
         );
  or02d0 U7936 ( .A1(n9875), .A2(n7429), .Z(n5155) );
  oai31d1 U7941 ( .B1(n11541), .B2(n11542), .B3(n6914), .A(n3937), .ZN(n11539)
         );
  oai21d1 U7943 ( .B1(n3939), .B2(n6914), .A(n5161), .ZN(n11543) );
  aoi31d1 U7955 ( .B1(n7666), .B2(n11546), .B3(n3910), .A(n7667), .ZN(n11542)
         );
  oai311d1 U7959 ( .C1(n11541), .C2(n11548), .C3(n7669), .A(n3953), .B(n6003), 
        .ZN(n11546) );
  oai21d1 U7960 ( .B1(n5178), .B2(n11549), .A(n8865), .ZN(n7669) );
  aoi31d1 U7968 ( .B1(n11550), .B2(n8090), .B3(n11551), .A(n6632), .ZN(n11548)
         );
  aoi22d1 U7976 ( .A1(n3957), .A2(n5769), .B1(n3957), .B2(n11553), .ZN(n11551)
         );
  oai211d1 U7977 ( .C1(n11554), .C2(n5187), .A(n4957), .B(n11550), .ZN(n11553)
         );
  aoi211d1 U7980 ( .C1(n5770), .C2(n7243), .A(n11557), .B(n11558), .ZN(n11554)
         );
  oan211d1 U7981 ( .C1(n6013), .C2(n6014), .B(n11559), .A(n6016), .ZN(n11558)
         );
  oai31d1 U7982 ( .B1(n11557), .B2(n11560), .B3(n11561), .A(n3824), .ZN(n11559) );
  aoi31d1 U7986 ( .B1(n3886), .B2(n5753), .B3(n11564), .A(n6022), .ZN(n11560)
         );
  aoi211d1 U7988 ( .C1(n3831), .C2(n11565), .A(n3829), .B(n11566), .ZN(n11564)
         );
  oan211d1 U7989 ( .C1(n11567), .C2(n6030), .B(n4698), .A(n6625), .ZN(n11566)
         );
  oan211d1 U7995 ( .C1(n11568), .C2(n11569), .B(n3879), .A(n11568), .ZN(n11567) );
  oai22d1 U7996 ( .A1(n11570), .A2(n3837), .B1(n3839), .B2(n10674), .ZN(n11569) );
  oai21d1 U7998 ( .B1(n7685), .B2(n11571), .A(images_bus[199]), .ZN(n6034) );
  aoim211d1 U8005 ( .C1(n5214), .C2(n11572), .A(n11573), .B(n11574), .ZN(
        n11570) );
  aoi31d1 U8006 ( .B1(n11572), .B2(n6040), .B3(n11575), .A(n4409), .ZN(n11574)
         );
  aoi22d1 U8011 ( .A1(n11578), .A2(n3853), .B1(n11579), .B2(n6046), .ZN(n11577) );
  oai211d1 U8017 ( .C1(n6050), .C2(n11580), .A(n3883), .B(n6052), .ZN(n11578)
         );
  aoi21d1 U8018 ( .B1(n5839), .B2(n3868), .A(n4314), .ZN(n6052) );
  aoi221d1 U8020 ( .B1(n11582), .B2(n6053), .C1(n3618), .C2(n6055), .A(n6057), 
        .ZN(n11580) );
  oai211d1 U8021 ( .C1(n11583), .C2(n5262), .A(n11257), .B(n5758), .ZN(n6057)
         );
  aoi321d1 U8025 ( .C1(n3862), .C2(n5275), .C3(n6062), .B1(n8082), .B2(n7708), 
        .A(n7710), .ZN(n11584) );
  oai21d1 U8026 ( .B1(images_bus[219]), .B2(n9929), .A(n11585), .ZN(n7710) );
  aon211d1 U8027 ( .C1(n9189), .C2(n11586), .B(n3619), .A(n3862), .ZN(n11585)
         );
  oai21d1 U8031 ( .B1(images_bus[225]), .B2(n3732), .A(images_bus[223]), .ZN(
        n5275) );
  aor22d1 U8046 ( .A1(n6062), .A2(n11587), .B1(n3721), .B2(n11588), .Z(n11582)
         );
  oai22d1 U8048 ( .A1(n11589), .A2(n6066), .B1(n11590), .B2(n3730), .ZN(n11587) );
  oan211d1 U8055 ( .C1(n11591), .C2(n5268), .B(n3742), .A(n11592), .ZN(n11590)
         );
  aoi31d1 U8059 ( .B1(n5274), .B2(n11593), .B3(n3672), .A(n5286), .ZN(n11591)
         );
  aon211d1 U8061 ( .C1(n3748), .C2(n11595), .B(n4691), .A(n6073), .ZN(n11593)
         );
  oai211d1 U8064 ( .C1(n11596), .C2(n9202), .A(n3753), .B(n3668), .ZN(n11595)
         );
  oai22d1 U8066 ( .A1(images_bus[231]), .A2(n9202), .B1(n6978), .B2(n11599), 
        .ZN(n6076) );
  oan211d1 U8072 ( .C1(n11600), .C2(n11601), .B(n3759), .A(n11602), .ZN(n11596) );
  aoi311d1 U8075 ( .C1(n3665), .C2(n6087), .C3(n11604), .A(n5301), .B(n10722), 
        .ZN(n11600) );
  oai21d1 U8076 ( .B1(n9626), .B2(n5300), .A(n6082), .ZN(n5301) );
  aoi21d1 U8077 ( .B1(n9207), .B2(images_bus[233]), .A(n6985), .ZN(n6082) );
  oan211d1 U8083 ( .C1(n11606), .C2(n5308), .B(n5309), .A(n5300), .ZN(n11604)
         );
  or02d0 U8084 ( .A1(n9949), .A2(n7413), .Z(n5300) );
  oan211d1 U8089 ( .C1(images_bus[239]), .C2(n6092), .B(n11608), .A(n10728), 
        .ZN(n11606) );
  aon211d1 U8090 ( .C1(n3800), .C2(n11609), .B(n11610), .A(n3773), .ZN(n11608)
         );
  oai211d1 U8096 ( .C1(n11611), .C2(n3779), .A(n6099), .B(n3775), .ZN(n11609)
         );
  oai21d1 U8098 ( .B1(n3778), .B2(n10735), .A(images_bus[241]), .ZN(n6095) );
  or02d0 U8099 ( .A1(n7729), .A2(n5544), .Z(n6099) );
  oai21d1 U8100 ( .B1(n11613), .B2(n5319), .A(n10407), .ZN(n7729) );
  aoi211d1 U8108 ( .C1(n6103), .C2(n11616), .A(n11617), .B(n6106), .ZN(n11611)
         );
  or02d0 U8109 ( .A1(n11610), .A2(n6105), .Z(n11617) );
  oai21d1 U8110 ( .B1(n10734), .B2(n7004), .A(images_bus[243]), .ZN(n6105) );
  or02d0 U8111 ( .A1(n9222), .A2(images_bus[245]), .Z(n7004) );
  oai211d1 U8112 ( .C1(n6108), .C2(n6109), .A(n2791), .B(n6110), .ZN(n11616)
         );
  aoim31d1 U8118 ( .B1(n11621), .B2(n7411), .B3(n6620), .A(n7742), .ZN(n11620)
         );
  oai21d1 U8123 ( .B1(n11622), .B2(n11623), .A(images_bus[251]), .ZN(n6620) );
  oai222d1 U8124 ( .A1(n11624), .A2(n8077), .B1(n11625), .B2(n7747), .C1(
        images_bus[253]), .C2(n11626), .ZN(n11621) );
  oai21d1 U8125 ( .B1(n3522), .B2(n9235), .A(n3790), .ZN(n7747) );
  aoi211d1 U8139 ( .C1(n5348), .C2(n6113), .A(n11627), .B(n11628), .ZN(n11624)
         );
  aoi31d1 U8140 ( .B1(n11629), .B2(images_bus[256]), .B3(n11630), .A(n4395), 
        .ZN(n11628) );
  oan211d1 U8143 ( .C1(n11632), .C2(n11633), .B(n3526), .A(n4435), .ZN(n11630)
         );
  aoi31d1 U8150 ( .B1(n3528), .B2(n8855), .B3(n11635), .A(n3568), .ZN(n11632)
         );
  aon211d1 U8152 ( .C1(images_bus[259]), .C2(n9240), .B(n8464), .A(n9239), 
        .ZN(n11636) );
  aoi22d1 U8159 ( .A1(n3529), .A2(n11638), .B1(n3530), .B2(n11633), .ZN(n11635) );
  aon211d1 U8160 ( .C1(n11639), .C2(n11640), .B(n4449), .A(n3510), .ZN(n11638)
         );
  aoi21d1 U8164 ( .B1(n3535), .B2(n11642), .A(n11643), .ZN(n11640) );
  aoi31d1 U8165 ( .B1(n3510), .B2(n4454), .B3(n11644), .A(n4456), .ZN(n11643)
         );
  aoi31d1 U8166 ( .B1(n3561), .B2(n11645), .B3(n3537), .A(n11646), .ZN(n11644)
         );
  aoi311d1 U8167 ( .C1(n3509), .C2(n4461), .C3(n11648), .A(n3541), .B(n4465), 
        .ZN(n11646) );
  aoi22d1 U8172 ( .A1(n4466), .A2(n11649), .B1(n4468), .B2(n11650), .ZN(n11648) );
  oai211d1 U8173 ( .C1(n3508), .C2(n3551), .A(n11652), .B(n4473), .ZN(n11650)
         );
  oai211d1 U8175 ( .C1(images_bus[285]), .C2(n3555), .A(n5414), .B(n11654), 
        .ZN(n8498) );
  aoi21d1 U8176 ( .B1(n3554), .B2(n6158), .A(n12169), .ZN(n11654) );
  oai31d1 U8179 ( .B1(n11655), .B2(n4475), .B3(n11649), .A(n4476), .ZN(n11652)
         );
  oai321d1 U8187 ( .C1(n4478), .C2(images_bus[289]), .C3(n5382), .B1(
        images_bus[287]), .B2(n9273), .A(n3494), .ZN(n4475) );
  oai22d1 U8189 ( .A1(n11656), .A2(n4478), .B1(n4479), .B2(n11657), .ZN(n11655) );
  aon211d1 U8190 ( .C1(n3473), .C2(n11658), .B(n4483), .A(n4484), .ZN(n11657)
         );
  oai31d1 U8192 ( .B1(n11661), .B2(n11662), .B3(n4488), .A(n3428), .ZN(n11660)
         );
  or02d0 U8196 ( .A1(n11663), .A2(n4675), .Z(n4488) );
  oan211d1 U8198 ( .C1(n7059), .C2(images_bus[295]), .B(n4677), .A(n5392), 
        .ZN(n11663) );
  aoi31d1 U8199 ( .B1(n3496), .B2(n4492), .B3(n11665), .A(n4495), .ZN(n11662)
         );
  aoi22d1 U8207 ( .A1(n11666), .A2(n3433), .B1(n4498), .B2(n11667), .ZN(n11665) );
  aoi21d1 U8211 ( .B1(n11669), .B2(n11670), .A(n4502), .ZN(n11666) );
  aon211d1 U8212 ( .C1(n3435), .C2(n11671), .B(n4505), .A(n3434), .ZN(n11670)
         );
  oai221d1 U8215 ( .B1(images_bus[304]), .B2(n11672), .C1(images_bus[305]), 
        .C2(n6181), .A(images_bus[303]), .ZN(n4505) );
  oai211d1 U8217 ( .C1(n11674), .C2(n4508), .A(n4509), .B(n11669), .ZN(n11671)
         );
  ora211d1 U8218 ( .C1(n7796), .C2(n11675), .A(images_bus[303]), .B(n11676), 
        .Z(n4509) );
  aoi31d1 U8220 ( .B1(n3456), .B2(n4307), .B3(n3457), .A(n11678), .ZN(n7789)
         );
  oan211d1 U8221 ( .C1(n11679), .C2(n7090), .B(images_bus[307]), .A(n5412), 
        .ZN(n11678) );
  aon211d1 U8223 ( .C1(n7797), .C2(n7395), .B(n7799), .A(n3457), .ZN(n11675)
         );
  oai21d1 U8225 ( .B1(n11680), .B2(n3450), .A(images_bus[311]), .ZN(n7799) );
  aoi21d1 U8227 ( .B1(n3449), .B2(n11680), .A(n9312), .ZN(n7797) );
  aoi31d1 U8243 ( .B1(n4518), .B2(n11684), .B3(n3495), .A(n7796), .ZN(n11682)
         );
  aor31d1 U8252 ( .B1(n4525), .B2(n11686), .B3(n11687), .A(n4517), .Z(n11684)
         );
  oai211d1 U8254 ( .C1(n4528), .C2(n4527), .A(n11688), .B(n4522), .ZN(n11686)
         );
  aon211d1 U8256 ( .C1(n3348), .C2(n4531), .B(n11691), .A(n4528), .ZN(n11688)
         );
  aoi311d1 U8262 ( .C1(n3346), .C2(n3368), .C3(n11695), .A(n4539), .B(n4538), 
        .ZN(n11692) );
  aoi221d1 U8266 ( .B1(n3371), .B2(n3347), .C1(n3413), .C2(n11700), .A(n4543), 
        .ZN(n11695) );
  oai21d1 U8267 ( .B1(images_bus[327]), .B2(n5438), .A(n6210), .ZN(n4543) );
  oai321d1 U8270 ( .C1(n11701), .C2(n7132), .C3(n3370), .B1(n11703), .B2(
        n10393), .A(n11704), .ZN(n11700) );
  oai21d1 U8272 ( .B1(n11706), .B2(n10393), .A(n4668), .ZN(n4554) );
  aoi221d1 U8274 ( .B1(n10071), .B2(n5726), .C1(n3410), .C2(n5633), .A(n11707), 
        .ZN(n11706) );
  oan211d1 U8275 ( .C1(n7132), .C2(n6230), .B(images_bus[331]), .A(n11708), 
        .ZN(n11707) );
  oaim21d1 U8290 ( .B1(n4558), .B2(n11711), .A(n11712), .ZN(n11701) );
  aoi221d1 U8292 ( .B1(n4559), .B2(n11714), .C1(n3379), .C2(n11715), .A(n4563), 
        .ZN(n11713) );
  oai211d1 U8296 ( .C1(n11717), .C2(n4565), .A(n4566), .B(n11718), .ZN(n11714)
         );
  aoi21d1 U8297 ( .B1(n3381), .B2(n11719), .A(n11715), .ZN(n11718) );
  aon211d1 U8299 ( .C1(n11720), .C2(n11721), .B(n11722), .A(n7135), .ZN(n7833)
         );
  aoi21d1 U8300 ( .B1(n3397), .B2(n11723), .A(n6258), .ZN(n11722) );
  oai211d1 U8302 ( .C1(images_bus[343]), .C2(n10081), .A(n11725), .B(
        images_bus[341]), .ZN(n11724) );
  oan211d1 U8318 ( .C1(n4981), .C2(n8575), .B(n3385), .A(n11728), .ZN(n7838)
         );
  aoi31d1 U8322 ( .B1(n3251), .B2(n11730), .B3(n11731), .A(n3386), .ZN(n11727)
         );
  aor31d1 U8326 ( .B1(n11731), .B2(n4577), .B3(n11732), .A(n4579), .Z(n11730)
         );
  aoi22d1 U8329 ( .A1(n3273), .A2(n11733), .B1(n4582), .B2(n11734), .ZN(n11732) );
  aon211d1 U8330 ( .C1(n11735), .C2(n11736), .B(n4586), .A(n3327), .ZN(n11734)
         );
  oan211d1 U8339 ( .C1(n11742), .C2(n11743), .B(n3320), .A(n3322), .ZN(n11735)
         );
  aoim211d1 U8349 ( .C1(n4599), .C2(n4598), .A(n3317), .B(n11745), .ZN(n11742)
         );
  oan211d1 U8350 ( .C1(n3279), .C2(n11746), .B(n11747), .A(n4597), .ZN(n11745)
         );
  nd13d1 U8351 ( .A1(n9388), .A2(n11748), .A3(n5480), .ZN(n4597) );
  oai211d1 U8353 ( .C1(n11749), .C2(n4607), .A(n11750), .B(n11751), .ZN(n11747) );
  aon211d1 U8355 ( .C1(n6316), .C2(n6318), .B(n7175), .A(n3313), .ZN(n11750)
         );
  aoi211d1 U8367 ( .C1(n3285), .C2(n11755), .A(n11756), .B(n6317), .ZN(n11749)
         );
  oai22d1 U8369 ( .A1(n11757), .A2(n4613), .B1(n11758), .B2(n4615), .ZN(n11756) );
  aoi311d1 U8370 ( .C1(n3293), .C2(n11759), .C3(n3290), .A(n11755), .B(n4620), 
        .ZN(n11758) );
  oai211d1 U8372 ( .C1(n8065), .C2(n8066), .A(n11760), .B(n11761), .ZN(n11759)
         );
  aoi211d1 U8373 ( .C1(n11762), .C2(n4624), .A(n3264), .B(n5043), .ZN(n11761)
         );
  aon211d1 U8376 ( .C1(n3309), .C2(n3307), .B(n8066), .A(n11765), .ZN(n4624)
         );
  oan211d1 U8380 ( .C1(n11767), .C2(n11768), .B(n3304), .A(n8067), .ZN(n11760)
         );
  oaim22d1 U8391 ( .A1(n11773), .A2(n8616), .B1(n11774), .B2(n3300), .ZN(
        n11767) );
  aoi311d1 U8399 ( .C1(n3294), .C2(n11775), .C3(n3165), .A(n4634), .B(n11774), 
        .ZN(n11773) );
  nd13d1 U8400 ( .A1(n8063), .A2(n8843), .A3(n11776), .ZN(n4634) );
  aoi21d1 U8401 ( .B1(n11777), .B2(n4969), .A(n11778), .ZN(n11776) );
  oan211d1 U8402 ( .C1(n3161), .C2(n7211), .B(images_bus[381]), .A(n8842), 
        .ZN(n11778) );
  aon211d1 U8403 ( .C1(n3163), .C2(n3168), .B(n8842), .A(n8845), .ZN(n11777)
         );
  oai211d1 U8420 ( .C1(n11781), .C2(n4638), .A(n3247), .B(n11782), .ZN(n11775)
         );
  oai31d1 U8422 ( .B1(n6365), .B2(images_bus[384]), .B3(n3248), .A(n11783), 
        .ZN(n5513) );
  aoi211d1 U8434 ( .C1(n3172), .C2(n11784), .A(n11785), .B(n11786), .ZN(n11781) );
  aoi31d1 U8435 ( .B1(n3149), .B2(n5528), .B3(n11788), .A(n10129), .ZN(n11786)
         );
  aoi22d1 U8440 ( .A1(n11790), .A2(n11791), .B1(n11792), .B2(n3181), .ZN(
        n11788) );
  oan211d1 U8442 ( .C1(n6379), .C2(n8634), .B(n11791), .A(n11794), .ZN(n5525)
         );
  aoi31d1 U8445 ( .B1(n11795), .B2(n5537), .B3(n11796), .A(n3183), .ZN(n11790)
         );
  aoi22d1 U8448 ( .A1(n11797), .A2(n5539), .B1(n3188), .B2(n11798), .ZN(n11796) );
  oai22d1 U8449 ( .A1(n5538), .A2(n3148), .B1(n11800), .B2(n3197), .ZN(n11798)
         );
  aoi221d1 U8451 ( .B1(n3202), .B2(n11801), .C1(n7902), .C2(n11802), .A(n5710), 
        .ZN(n11800) );
  oai21d1 U8452 ( .B1(n5910), .B2(n3205), .A(n7899), .ZN(n5710) );
  oai22d1 U8457 ( .A1(n11219), .A2(n7898), .B1(n11806), .B2(n9437), .ZN(n7902)
         );
  oai221d1 U8460 ( .B1(n11807), .B2(n8059), .C1(n11808), .C2(n7900), .A(n3210), 
        .ZN(n11801) );
  oai21d1 U8462 ( .B1(n11219), .B2(images_bus[403]), .A(n11810), .ZN(n11809)
         );
  oai21d1 U8465 ( .B1(n6409), .B2(n6416), .A(n11219), .ZN(n7900) );
  aoi211d1 U8474 ( .C1(n5562), .C2(n11802), .A(n11811), .B(n5559), .ZN(n11807)
         );
  oai21d1 U8475 ( .B1(n3231), .B2(n4961), .A(n4685), .ZN(n5559) );
  aoi21d1 U8476 ( .B1(n5709), .B2(n5554), .A(n11812), .ZN(n4685) );
  oai221d1 U8479 ( .B1(n8058), .B2(n3147), .C1(n11814), .C2(n8057), .A(n7907), 
        .ZN(n11811) );
  aoi221d1 U8481 ( .B1(n11815), .B2(n5556), .C1(n11003), .C2(n11816), .A(n5557), .ZN(n11814) );
  oan211d1 U8483 ( .C1(n4900), .C2(n5709), .B(n11009), .A(n11818), .ZN(n4694)
         );
  oai22d1 U8486 ( .A1(n4901), .A2(n3027), .B1(n11819), .B2(n4704), .ZN(n11816)
         );
  aoi211d1 U8487 ( .C1(n3034), .C2(n11820), .A(n5707), .B(n4705), .ZN(n11819)
         );
  oai22d1 U8488 ( .A1(images_bus[413]), .A2(n3035), .B1(n7915), .B2(n11821), 
        .ZN(n4705) );
  oai21d1 U8491 ( .B1(n5706), .B2(n4702), .A(n11822), .ZN(n5707) );
  aon211d1 U8492 ( .C1(n4710), .C2(n4955), .B(n3039), .A(n3034), .ZN(n11822)
         );
  oai22d1 U8499 ( .A1(n3041), .A2(n4956), .B1(n11824), .B2(n4707), .ZN(n11820)
         );
  aoi221d1 U8501 ( .B1(n4955), .B2(n3047), .C1(n4715), .C2(n11825), .A(n7268), 
        .ZN(n11824) );
  oai21d1 U8502 ( .B1(n5237), .B2(n4720), .A(n3048), .ZN(n7268) );
  oai221d1 U8508 ( .B1(n11826), .B2(n3057), .C1(n4646), .C2(n4724), .A(n7272), 
        .ZN(n11825) );
  aoi221d1 U8509 ( .B1(n5584), .B2(n3056), .C1(n7366), .C2(n4729), .A(n4952), 
        .ZN(n7272) );
  oai21d1 U8510 ( .B1(images_bus[421]), .B2(n3127), .A(n11827), .ZN(n4952) );
  oai21d1 U8514 ( .B1(n4730), .B2(n4731), .A(n4734), .ZN(n5584) );
  aoi21d1 U8515 ( .B1(n5980), .B2(n7935), .A(n11829), .ZN(n4734) );
  aoi221d1 U8541 ( .B1(n3064), .B2(n11831), .C1(n8694), .C2(n6465), .A(n5587), 
        .ZN(n11826) );
  oai21d1 U8542 ( .B1(n5140), .B2(n5589), .A(n7364), .ZN(n5587) );
  oai221d1 U8546 ( .B1(n11832), .B2(n5597), .C1(n5140), .C2(n3073), .A(n3070), 
        .ZN(n11831) );
  oai21d1 U8548 ( .B1(n4411), .B2(n5703), .A(n5593), .ZN(n9472) );
  aoi221d1 U8566 ( .B1(n7287), .B2(n11834), .C1(n4749), .C2(n5702), .A(n7284), 
        .ZN(n11832) );
  oai31d1 U8567 ( .B1(n10382), .B2(n5495), .B3(n3086), .A(n3080), .ZN(n7284)
         );
  oai221d1 U8569 ( .B1(n7962), .B2(n10382), .C1(n4411), .C2(n3120), .A(n5606), 
        .ZN(n11835) );
  oai22d1 U8570 ( .A1(n3120), .A2(n5902), .B1(n11836), .B2(n5600), .ZN(n5606)
         );
  aoi21d1 U8575 ( .B1(n5494), .B2(n7963), .A(n11837), .ZN(n7962) );
  aor21d1 U8583 ( .B1(n7963), .B2(n3117), .A(n7957), .Z(n4749) );
  oai211d1 U8586 ( .C1(n3090), .C2(n4945), .A(n5608), .B(n11841), .ZN(n11834)
         );
  aoi311d1 U8587 ( .C1(n7976), .C2(n6554), .C3(n3088), .A(n11843), .B(n11844), 
        .ZN(n11841) );
  aoi211d1 U8588 ( .C1(n11845), .C2(n7975), .A(n4763), .B(n9490), .ZN(n11844)
         );
  aoi22d1 U8590 ( .A1(n4778), .A2(n4894), .B1(n8736), .B2(n6500), .ZN(n7975)
         );
  aoi22d1 U8593 ( .A1(n3016), .A2(n11846), .B1(n4777), .B2(n7974), .ZN(n11845)
         );
  oai211d1 U8598 ( .C1(n11847), .C2(n5635), .A(n5628), .B(n11848), .ZN(n11846)
         );
  aoi21d1 U8599 ( .B1(n6503), .B2(n4942), .A(n4781), .ZN(n11848) );
  aor21d1 U8600 ( .B1(n4779), .B2(n7972), .A(n5627), .Z(n4781) );
  oaim21d1 U8602 ( .B1(n4788), .B2(n2925), .A(n4785), .ZN(n6503) );
  oai21d1 U8606 ( .B1(n8039), .B2(n11850), .A(n11851), .ZN(n4790) );
  oai211d1 U8607 ( .C1(n11852), .C2(n8031), .A(n5727), .B(n2938), .ZN(n11851)
         );
  aoi211d1 U8628 ( .C1(n4791), .C2(n4942), .A(n11855), .B(n2942), .ZN(n11847)
         );
  aoi21d1 U8630 ( .B1(n4802), .B2(n2944), .A(n4797), .ZN(n5637) );
  aon211d1 U8631 ( .C1(n8039), .C2(images_bus[451]), .B(n3007), .A(n11856), 
        .ZN(n4797) );
  oai221d1 U8634 ( .B1(n9510), .B2(n11858), .C1(images_bus[453]), .C2(n3005), 
        .A(n11859), .ZN(n4802) );
  oai22d1 U8636 ( .A1(n5639), .A2(n11861), .B1(n11862), .B2(n5641), .ZN(n11855) );
  aoim211d1 U8639 ( .C1(n11861), .C2(n2955), .A(n11863), .B(n2952), .ZN(n11862) );
  aoi21d1 U8641 ( .B1(n4812), .B2(n2953), .A(n4809), .ZN(n6515) );
  oai22d1 U8642 ( .A1(n2955), .A2(n7360), .B1(n8756), .B2(n11864), .ZN(n4809)
         );
  oai22d1 U8645 ( .A1(n5129), .A2(n4815), .B1(n7316), .B2(n11866), .ZN(n4812)
         );
  oai22d1 U8648 ( .A1(n11867), .A2(n4807), .B1(n11868), .B2(n2954), .ZN(n11863) );
  oai22d1 U8650 ( .A1(n4804), .A2(n4803), .B1(n4815), .B2(n4807), .ZN(n6517)
         );
  aoi211d1 U8653 ( .C1(n2991), .C2(n11869), .A(n11870), .B(n5651), .ZN(n11867)
         );
  aoim2m11d1 U8655 ( .C1(images_bus[463]), .C2(n11871), .B(n11872), .A(n8760), 
        .ZN(n4817) );
  aoi22d1 U8657 ( .A1(n7982), .A2(n2990), .B1(n7359), .B2(n8759), .ZN(n11872)
         );
  aoi22d1 U8659 ( .A1(n2994), .A2(n9525), .B1(n2990), .B2(n11873), .ZN(n11871)
         );
  oai22d1 U8660 ( .A1(n11868), .A2(n2997), .B1(n11874), .B2(n5654), .ZN(n11870) );
  aoi211d1 U8663 ( .C1(n2961), .C2(n11869), .A(n11875), .B(n5657), .ZN(n11874)
         );
  aon211d1 U8664 ( .C1(n4828), .C2(n4937), .B(n7357), .A(n11876), .ZN(n5657)
         );
  aoi21d1 U8670 ( .B1(n2986), .B2(n4820), .A(n7986), .ZN(n4828) );
  oaim21d1 U8671 ( .B1(n2986), .B2(n11878), .A(n11879), .ZN(n7986) );
  aon211d1 U8672 ( .C1(n4838), .C2(n11880), .B(n11881), .A(n2968), .ZN(n11879)
         );
  oai22d1 U8674 ( .A1(n11883), .A2(n5659), .B1(n11884), .B2(n5661), .ZN(n11875) );
  aoi211d1 U8676 ( .C1(n5662), .C2(n11885), .A(n11886), .B(n2972), .ZN(n11884)
         );
  oaim21d1 U8679 ( .B1(n7992), .B2(n4933), .A(n7990), .ZN(n4842) );
  oan211d1 U8680 ( .C1(n11880), .C2(n5798), .B(n4840), .A(n11887), .ZN(n7990)
         );
  oai21d1 U8682 ( .B1(images_bus[473]), .B2(n2979), .A(n11888), .ZN(n7992) );
  oai22d1 U8685 ( .A1(n5666), .A2(n11883), .B1(n11889), .B2(n5668), .ZN(n11886) );
  aoi221d1 U8687 ( .B1(n2978), .B2(n11890), .C1(n5671), .C2(n11885), .A(n5672), 
        .ZN(n11889) );
  oai21d1 U8688 ( .B1(n2825), .B2(n6542), .A(n2818), .ZN(n5672) );
  oai22d1 U8690 ( .A1(n8782), .A2(n4934), .B1(n6542), .B2(n8792), .ZN(n4935)
         );
  oai221d1 U8694 ( .B1(n6079), .B2(n4931), .C1(n2829), .C2(n11893), .A(n11894), 
        .ZN(n11891) );
  oai21d1 U8698 ( .B1(n2829), .B2(n6542), .A(n4934), .ZN(n5671) );
  or02d0 U8699 ( .A1(n7356), .A2(n7331), .Z(n4934) );
  oai22d1 U8700 ( .A1(n11895), .A2(n4929), .B1(n5675), .B2(n11896), .ZN(n11890) );
  aoi321d1 U8711 ( .C1(n2851), .C2(n11899), .C3(n5678), .B1(n5679), .B2(n11900), .A(n11901), .ZN(n11895) );
  oai21d1 U8712 ( .B1(n4930), .B2(n11896), .A(n5682), .ZN(n11901) );
  aoi21d1 U8713 ( .B1(n7349), .B2(n5679), .A(n2843), .ZN(n5682) );
  aon211d1 U8715 ( .C1(n11903), .C2(n7337), .B(n7338), .A(n5678), .ZN(n6546)
         );
  oai21d1 U8716 ( .B1(images_bus[481]), .B2(n2913), .A(n11904), .ZN(n7338) );
  oai21d1 U8718 ( .B1(n4869), .B2(images_bus[483]), .A(n9555), .ZN(n7349) );
  aoi21d1 U8720 ( .B1(n7337), .B2(n5678), .A(n2844), .ZN(n4930) );
  oai211d1 U8721 ( .C1(n2836), .C2(n4870), .A(n2853), .B(n11908), .ZN(n11900)
         );
  aoi22d1 U8722 ( .A1(n2855), .A2(n11909), .B1(n2856), .B2(n11910), .ZN(n11908) );
  oai211d1 U8723 ( .C1(n2835), .C2(n2870), .A(n2867), .B(n11912), .ZN(n11910)
         );
  aoi22d1 U8724 ( .A1(n2869), .A2(n11913), .B1(n4878), .B2(n11914), .ZN(n11912) );
  oai211d1 U8726 ( .C1(n11915), .C2(n4884), .A(n4885), .B(n11916), .ZN(n11913)
         );
  aoi21d1 U8727 ( .B1(n4879), .B2(n11914), .A(n2873), .ZN(n11916) );
  aoi221d1 U8729 ( .B1(n2880), .B2(n11918), .C1(n8815), .C2(n11919), .A(n8809), 
        .ZN(n7352) );
  oai221d1 U8730 ( .B1(n5124), .B2(n11921), .C1(images_bus[491]), .C2(n2911), 
        .A(n11923), .ZN(n8809) );
  oan211d1 U8734 ( .C1(n4924), .C2(n4393), .B(n11186), .A(n11925), .ZN(n11924)
         );
  nd13d1 U8737 ( .A1(n11919), .A2(n11921), .A3(n11927), .ZN(n4879) );
  aoi21d1 U8738 ( .B1(n11918), .B2(n11186), .A(n8828), .ZN(n11927) );
  oai21d1 U8739 ( .B1(n11142), .B2(n11928), .A(n2911), .ZN(n11921) );
  aoi211d1 U8760 ( .C1(n11933), .C2(n4920), .A(n11934), .B(n4921), .ZN(n11915)
         );
  oaim21d1 U8761 ( .B1(n2884), .B2(n8013), .A(n8009), .ZN(n4921) );
  oai22d1 U8767 ( .A1(n11935), .A2(n2883), .B1(n11936), .B2(n8008), .ZN(n11934) );
  aoi221d1 U8769 ( .B1(n2833), .B2(n2907), .C1(n2905), .C2(n11939), .A(n11940), 
        .ZN(n11936) );
  oai211d1 U8770 ( .C1(n2834), .C2(n4891), .A(n11942), .B(n8014), .ZN(n11940)
         );
  aon211d1 U8771 ( .C1(n2891), .C2(n12173), .B(n11943), .A(n2903), .ZN(n8014)
         );
  oai211d1 U8773 ( .C1(n4909), .C2(n11944), .A(n4898), .B(n2903), .ZN(n11942)
         );
  oaim22d1 U8774 ( .A1(n11945), .A2(n4904), .B1(n4908), .B2(n11939), .ZN(
        n11944) );
  oan211d1 U8775 ( .C1(n4916), .C2(n11939), .B(n8827), .A(n11946), .ZN(n11945)
         );
  aoi31d1 U8776 ( .B1(n8826), .B2(n8024), .B3(n11947), .A(n10339), .ZN(n11946)
         );
  oan211d1 U8778 ( .C1(n8020), .C2(n11948), .B(n8021), .A(n11949), .ZN(n11947)
         );
  oai21d1 U8780 ( .B1(n11951), .B2(n2899), .A(n11952), .ZN(n8021) );
  nd13d1 U8782 ( .A1(n4916), .A2(n4914), .A3(n2834), .ZN(n11948) );
  oai211d1 U8786 ( .C1(n10341), .C2(n2809), .A(n11181), .B(n2900), .ZN(n8826)
         );
  aoi31d1 U8802 ( .B1(N15554), .B2(n11953), .B3(n2896), .A(n11954), .ZN(n8827)
         );
  aor21d1 U8807 ( .B1(n9579), .B2(n4908), .A(n11956), .Z(n4909) );
  oan211d1 U8808 ( .C1(n2894), .C2(images_bus[503]), .B(n8823), .A(n4904), 
        .ZN(n11956) );
  or03d0 U8867 ( .A1(n11914), .A2(n8815), .A3(n11959), .Z(n11933) );
  oaim21d1 U8882 ( .B1(n11960), .B2(n4872), .A(n8803), .ZN(n4874) );
  oai21d1 U8901 ( .B1(n11962), .B2(n8801), .A(n8802), .ZN(n11961) );
  aon211d1 U8903 ( .C1(images_bus[484]), .C2(images_bus[483]), .B(n4870), .A(
        n11963), .ZN(n7350) );
  aon211d1 U8904 ( .C1(n11962), .C2(n11960), .B(n11964), .A(n8802), .ZN(n11963) );
  oai21d1 U8917 ( .B1(n11194), .B2(n2863), .A(n4869), .ZN(n4870) );
  aoim21d1 U8944 ( .B1(n4869), .B2(n7344), .A(n4860), .ZN(n7346) );
  aoi21d1 U8977 ( .B1(n4840), .B2(n7987), .A(n4839), .ZN(n5666) );
  aon211d1 U9002 ( .C1(n2968), .C2(n4838), .B(n4830), .A(n2962), .ZN(n5659) );
  aoi21d1 U9024 ( .B1(n2986), .B2(n2962), .A(n4821), .ZN(n6528) );
  aoi21d1 U9025 ( .B1(n11971), .B2(n2966), .A(n11873), .ZN(n4821) );
  oai21d1 U9043 ( .B1(n2998), .B2(n2999), .A(n4814), .ZN(n6527) );
  oai22d1 U9061 ( .A1(n2992), .A2(n7358), .B1(n11972), .B2(n7359), .ZN(n4822)
         );
  aoi22d1 U9103 ( .A1(n2941), .A2(n3007), .B1(n4800), .B2(n2944), .ZN(n5639)
         );
  oan211d1 U9150 ( .C1(n3109), .C2(n4763), .B(n4761), .A(n4301), .ZN(n11843)
         );
  oai21d1 U9158 ( .B1(n3103), .B2(n3099), .A(n4943), .ZN(n7976) );
  aoi21d1 U9167 ( .B1(n4772), .B2(n3089), .A(n3091), .ZN(n5608) );
  oai321d1 U9172 ( .C1(n6487), .C2(images_bus[439]), .C3(n3110), .B1(n6561), 
        .B2(n8053), .A(n11976), .ZN(n4772) );
  aon211d1 U9173 ( .C1(n11071), .C2(n12167), .B(n11977), .A(n4764), .ZN(n11976) );
  aoi21d1 U9180 ( .B1(n11071), .B2(n4764), .A(n6485), .ZN(n8053) );
  oai22d1 U9293 ( .A1(n3030), .A2(n11009), .B1(n3035), .B2(n4704), .ZN(n4696)
         );
  oai21d1 U9308 ( .B1(n3227), .B2(n3214), .A(n6583), .ZN(n5556) );
  aoi21d1 U9323 ( .B1(n5552), .B2(n3231), .A(n5554), .ZN(n8058) );
  aoi21d1 U9364 ( .B1(n9437), .B2(n5529), .A(n4671), .ZN(n5538) );
  oai21d1 U9369 ( .B1(n3194), .B2(n4667), .A(n3190), .ZN(n5539) );
  aon211d1 U9376 ( .C1(n11985), .C2(n4963), .B(n4673), .A(n3188), .ZN(n11986)
         );
  aoim211d1 U9411 ( .C1(n11990), .C2(n3242), .A(n4659), .B(n5982), .ZN(n5528)
         );
  aoi21d1 U9420 ( .B1(n8634), .B2(n6591), .A(n3182), .ZN(n11990) );
  aoim31d1 U9422 ( .B1(n6380), .B2(images_bus[395]), .B3(n6379), .A(n5625), 
        .ZN(n4660) );
  aoi211d1 U9439 ( .C1(n3173), .C2(n4652), .A(n4642), .B(n11994), .ZN(n5515)
         );
  oan211d1 U9440 ( .C1(n4648), .C2(n3175), .B(n3170), .A(n4645), .ZN(n11994)
         );
  aoi221d1 U9514 ( .B1(n5818), .B2(n10953), .C1(n9606), .C2(n11766), .A(n4304), 
        .ZN(n8065) );
  or02d0 U9547 ( .A1(n11746), .A2(n4423), .Z(n11755) );
  oan211d1 U9577 ( .C1(n7385), .C2(n11999), .B(n5997), .A(n9388), .ZN(n4599)
         );
  aoim31d1 U9586 ( .B1(n7169), .B2(n11752), .B3(n7381), .A(n12165), .ZN(n11748) );
  aoi321d1 U9609 ( .C1(n3273), .C2(n5732), .C3(n3330), .B1(n4979), .B2(n4582), 
        .A(n8072), .ZN(n4577) );
  oai22d1 U9645 ( .A1(n6277), .A2(n9374), .B1(images_bus[349]), .B2(n6275), 
        .ZN(n7845) );
  oai22d1 U9681 ( .A1(n6243), .A2(n9354), .B1(n3378), .B2(n12006), .ZN(n7831)
         );
  oai211d1 U9713 ( .C1(n4427), .C2(n12011), .A(n3404), .B(n12012), .ZN(n4558)
         );
  aon211d1 U9716 ( .C1(n6602), .C2(n6237), .B(n9346), .A(n12013), .ZN(n12011)
         );
  oai21d1 U9770 ( .B1(n3366), .B2(n5737), .A(n3419), .ZN(n4531) );
  aoi211d1 U9806 ( .C1(n4992), .C2(n7804), .A(n7807), .B(n12020), .ZN(n4518)
         );
  aoi321d1 U9848 ( .C1(n12022), .C2(n5164), .C3(n10825), .B1(n3465), .B2(n5636), .A(n12023), .ZN(n12021) );
  oan211d1 U9849 ( .C1(n12024), .C2(n10828), .B(n8524), .A(n4502), .ZN(n12023)
         );
  aoi31d1 U9856 ( .B1(n3460), .B2(n6183), .B3(n11668), .A(n4436), .ZN(n12024)
         );
  oai21d1 U9888 ( .B1(n4997), .B2(n11661), .A(n3472), .ZN(n11659) );
  aoi322d1 U9943 ( .C1(n3545), .C2(n5834), .C3(n3543), .A1(n9255), .A2(n12030), 
        .B1(n4468), .B2(n8497), .ZN(n12028) );
  oai21d1 U9944 ( .B1(n12031), .B2(n6151), .A(images_bus[281]), .ZN(n8497) );
  aoi21d1 U9946 ( .B1(n3553), .B2(n12026), .A(n12033), .ZN(n12031) );
  aoi211d1 U9975 ( .C1(n3558), .C2(n4311), .A(n5742), .B(n9620), .ZN(n12027)
         );
  aoim211d1 U9985 ( .C1(n12035), .C2(n6616), .A(n7152), .B(n8482), .ZN(n4454)
         );
  aoi21d1 U9988 ( .B1(n3560), .B2(n7766), .A(n5933), .ZN(n12035) );
  aon211d1 U9990 ( .C1(n3540), .C2(n5060), .B(n9620), .A(n9998), .ZN(n12036)
         );
  nd13d1 U10024 ( .A1(n11633), .A2(n6134), .A3(n8855), .ZN(n12038) );
  oai21d1 U10049 ( .B1(n6128), .B2(n12044), .A(n12045), .ZN(n12043) );
  aon211d1 U10050 ( .C1(n8471), .C2(n12042), .B(n6388), .A(n3530), .ZN(n12045)
         );
  aon211d1 U10051 ( .C1(n3533), .C2(n5644), .B(n7152), .A(n3532), .ZN(n12044)
         );
  aoi21d1 U10102 ( .B1(n7411), .B2(n3784), .A(n7740), .ZN(n6108) );
  oai21d1 U10119 ( .B1(n7003), .B2(n10734), .A(n5328), .ZN(n6103) );
  or02d0 U10147 ( .A1(n10726), .A2(images_bus[237]), .Z(n5303) );
  aoi21d1 U10220 ( .B1(n7704), .B2(n3866), .A(n3867), .ZN(n6050) );
  oai21d1 U10227 ( .B1(n5248), .B2(n6961), .A(n5240), .ZN(n12052) );
  oan211d1 U10241 ( .C1(n8084), .C2(n5761), .B(n5219), .A(n8404), .ZN(n6040)
         );
  oai211d1 U10242 ( .C1(images_bus[205]), .C2(n11259), .A(images_bus[203]), 
        .B(images_bus[204]), .ZN(n8404) );
  oai21d1 U10246 ( .B1(images_bus[207]), .B2(n5227), .A(n4462), .ZN(n5761) );
  oai321d1 U10250 ( .C1(n5227), .C2(n3876), .C3(n5225), .B1(n3848), .B2(n12054), .A(n12055), .ZN(n8084) );
  aon211d1 U10251 ( .C1(n3871), .C2(n3854), .B(n5068), .A(n7691), .ZN(n12055)
         );
  aon211d1 U10268 ( .C1(n3875), .C2(n5234), .B(n5548), .A(n3874), .ZN(n12054)
         );
  or02d0 U10285 ( .A1(n11568), .A2(n5210), .Z(n11573) );
  oai21d1 U10287 ( .B1(images_bus[203]), .B2(n6943), .A(images_bus[201]), .ZN(
        n8400) );
  aoim21d1 U10340 ( .B1(n4958), .B2(n8380), .A(n9147), .ZN(n8090) );
  oai22d1 U10341 ( .A1(n12059), .A2(n3958), .B1(n12061), .B2(n12060), .ZN(
        n9147) );
  aoi221d1 U10371 ( .B1(n5774), .B2(n3945), .C1(n11552), .C2(n6003), .A(n4316), 
        .ZN(n7666) );
  nd13d1 U10551 ( .A1(n11462), .A2(n6651), .A3(images_bus[119]), .ZN(n11468)
         );
  aoim21d1 U10572 ( .B1(n11470), .B2(n6829), .A(n5447), .ZN(n7600) );
  oai21d1 U10665 ( .B1(images_bus[97]), .B2(n5031), .A(images_bus[95]), .ZN(
        n5878) );
  aoi321d1 U10690 ( .C1(n4170), .C2(n4061), .C3(n8104), .B1(n4973), .B2(n4168), 
        .A(n7447), .ZN(n7564) );
  aoi21d1 U10733 ( .B1(n5958), .B2(n4178), .A(n11407), .ZN(n5840) );
  aon211d1 U10757 ( .C1(n5828), .C2(n5691), .B(n7182), .A(n5821), .ZN(n8244)
         );
  nd13d1 U10759 ( .A1(n6748), .A2(n4184), .A3(N8868), .ZN(n6750) );
  oai22d1 U10850 ( .A1(n4248), .A2(n10493), .B1(images_bus[45]), .B2(n5800), 
        .ZN(n6706) );
  aoi21d1 U10881 ( .B1(n4754), .B2(n4233), .A(n4243), .ZN(n6687) );
  aon211d1 U10905 ( .C1(n4227), .C2(n8176), .B(n8125), .A(n7487), .ZN(n11334)
         );
  aoi21d1 U10979 ( .B1(n5315), .B2(n5794), .A(n6975), .ZN(n9645) );
  nd04d1 U3 ( .A1(n3578), .A2(n3579), .A3(n3580), .A4(n3581), .ZN(n12093) );
  nd04d1 U1064 ( .A1(n3607), .A2(n3608), .A3(n3609), .A4(n3610), .ZN(n12101)
         );
  nr03d1 U1077 ( .A1(n3617), .A2(n2783), .A3(n2777), .ZN(n3593) );
  an02d1 U1116 ( .A1(n3646), .A2(n2754), .Z(n3585) );
  an03d1 U1123 ( .A1(n3647), .A2(n2770), .A3(n3652), .Z(n3584) );
  an02d1 U1127 ( .A1(n493), .A2(n658), .Z(n3647) );
  nr03d1 U1130 ( .A1(n3652), .A2(n3651), .A3(n3655), .ZN(n3648) );
  nd04d1 U1156 ( .A1(n3656), .A2(n2775), .A3(n2777), .A4(n3654), .ZN(n3682) );
  nd04d1 U1164 ( .A1(n2770), .A2(reading_compare), .A3(n493), .A4(n2781), .ZN(
        n3686) );
  nr03d1 U1169 ( .A1(n3676), .A2(N5285), .A3(n3657), .ZN(n3649) );
  nd04d1 U1179 ( .A1(n3693), .A2(n3694), .A3(n3695), .A4(n3696), .ZN(n3691) );
  nd04d1 U1186 ( .A1(n3701), .A2(n2759), .A3(n3702), .A4(n3703), .ZN(n3690) );
  nr03d1 U1187 ( .A1(n3704), .A2(n6), .A3(n3705), .ZN(n3703) );
  nr04d1 U1205 ( .A1(compare_in_progress), .A2(hashes_ready), .A3(
        reading_compare), .A4(reading_current), .ZN(n3588) );
  nr03d1 U1781 ( .A1(N3232), .A2(N3233), .A3(N3231), .ZN(n4193) );
  nr03d1 U1787 ( .A1(n12210), .A2(N3231), .A3(n12211), .ZN(n4198) );
  nr03d1 U1790 ( .A1(n12210), .A2(N3232), .A3(n12212), .ZN(n4200) );
  nr03d1 U1793 ( .A1(N3231), .A2(N3232), .A3(n12210), .ZN(n4202) );
  nr03d1 U1796 ( .A1(n12211), .A2(N3233), .A3(n12212), .ZN(n4204) );
  nr03d1 U1799 ( .A1(N3231), .A2(N3233), .A3(n12211), .ZN(n4206) );
  nr03d1 U1806 ( .A1(N3232), .A2(N3233), .A3(n12212), .ZN(n4208) );
  nr03d1 U1811 ( .A1(n12211), .A2(n12210), .A3(n12212), .ZN(n4211) );
  nr03d1 U1827 ( .A1(n4237), .A2(new_reference_is_done), .A3(n2778), .ZN(n4236) );
  an02d1 U2274 ( .A1(n4362), .A2(N3878), .Z(n4329) );
  an02d1 U2477 ( .A1(n4362), .A2(n2789), .Z(n4345) );
  nd12d1 U2492 ( .A1(n4237), .A2(n4235), .ZN(n4375) );
  an02d1 U2493 ( .A1(n2771), .A2(N4760), .Z(n4235) );
  nr04d1 U2779 ( .A1(count_image[1]), .A2(count_image[0]), .A3(\lt_82/A[5] ), 
        .A4(\lt_82/A[4] ), .ZN(n4378) );
  nr03d1 U2782 ( .A1(count_image[6]), .A2(count_image[8]), .A3(count_image[7]), 
        .ZN(n4377) );
  an03d1 U2787 ( .A1(n2788), .A2(n2789), .A3(N3855), .Z(n4355) );
  nr04d1 U2790 ( .A1(n4379), .A2(n4380), .A3(n4381), .A4(n4382), .ZN(N26366)
         );
  nd04d1 U2791 ( .A1(n3856), .A2(n3795), .A3(n4385), .A4(n4386), .ZN(n4382) );
  nr04d1 U2792 ( .A1(n4387), .A2(n4388), .A3(n4389), .A4(n4390), .ZN(n4386) );
  nr03d1 U2794 ( .A1(n3781), .A2(n4394), .A3(n4395), .ZN(n4385) );
  nd04d1 U2795 ( .A1(n3792), .A2(n3574), .A3(n4398), .A4(n4399), .ZN(n4381) );
  nr04d1 U2796 ( .A1(n4400), .A2(n4401), .A3(n4402), .A4(n4403), .ZN(n4399) );
  nr03d1 U2798 ( .A1(n4407), .A2(n4016), .A3(n4409), .ZN(n4398) );
  nd04d1 U2800 ( .A1(n3725), .A2(n4412), .A3(n4413), .A4(n4414), .ZN(n4380) );
  nr04d1 U2801 ( .A1(n4415), .A2(n3934), .A3(n4417), .A4(n4418), .ZN(n4414) );
  nr03d1 U2803 ( .A1(n4422), .A2(n4023), .A3(n4424), .ZN(n4413) );
  nd04d1 U2805 ( .A1(n3805), .A2(n3862), .A3(n4428), .A4(n4429), .ZN(n4379) );
  nr04d1 U2806 ( .A1(n4430), .A2(n4431), .A3(n4432), .A4(n4433), .ZN(n4429) );
  nd04d1 U2820 ( .A1(n4477), .A2(n4485), .A3(n4486), .A4(n4487), .ZN(n4482) );
  nr04d1 U2836 ( .A1(n4533), .A2(n4534), .A3(n4535), .A4(n4536), .ZN(n4532) );
  nr04d1 U2838 ( .A1(n4541), .A2(n4542), .A3(n4543), .A4(n4538), .ZN(n4540) );
  nr04d1 U2847 ( .A1(n4570), .A2(n4571), .A3(n4569), .A4(n3384), .ZN(n4564) );
  nr04d1 U2858 ( .A1(n4609), .A2(n4610), .A3(n4611), .A4(n4605), .ZN(n4606) );
  nr04d1 U2866 ( .A1(n4641), .A2(n4642), .A3(n4643), .A4(n4644), .ZN(n4637) );
  nr03d1 U2950 ( .A1(n7050), .A2(n4924), .A3(n5894), .ZN(n4923) );
  nd12d1 U2951 ( .A1(n4867), .A2(n4925), .ZN(n4877) );
  nd12d1 U2961 ( .A1(n4831), .A2(n4936), .ZN(n4849) );
  an02d1 U2966 ( .A1(n4940), .A2(n2933), .Z(n4805) );
  an03d1 U2972 ( .A1(n4753), .A2(n4945), .A3(n4301), .Z(n4760) );
  an03d1 U2986 ( .A1(n4674), .A2(n4961), .A3(n5518), .Z(n4684) );
  nr03d1 U2995 ( .A1(n4969), .A2(n4970), .A3(n4632), .ZN(n4639) );
  an02d1 U3000 ( .A1(n4975), .A2(n4616), .Z(n4612) );
  nr03d1 U3003 ( .A1(n4581), .A2(n4978), .A3(n4979), .ZN(n4594) );
  nr03d1 U3005 ( .A1(n4569), .A2(n4981), .A3(n4982), .ZN(n4573) );
  nd12d1 U3006 ( .A1(n4562), .A2(n4983), .ZN(n4569) );
  an03d1 U3008 ( .A1(n4986), .A2(n4557), .A3(n4987), .Z(n4555) );
  an02d1 U3009 ( .A1(n4546), .A2(n4988), .Z(n4557) );
  nr03d1 U3010 ( .A1(n4989), .A2(n4541), .A3(n4990), .ZN(n4546) );
  nr03d1 U3014 ( .A1(n4519), .A2(n4992), .A3(n4993), .ZN(n4529) );
  an03d1 U3021 ( .A1(n5000), .A2(images_bus[288]), .A3(n4310), .Z(n4477) );
  nd12d1 U3025 ( .A1(n4452), .A2(n5002), .ZN(n4458) );
  nr03d1 U3028 ( .A1(n5006), .A2(n5007), .A3(n5008), .ZN(n4428) );
  nd04d1 U3030 ( .A1(n5010), .A2(n5011), .A3(n5012), .A4(n5013), .ZN(n4432) );
  nr04d1 U3031 ( .A1(n5014), .A2(n5015), .A3(n5016), .A4(n5017), .ZN(n5013) );
  an04d1 U3033 ( .A1(n5022), .A2(n5023), .A3(n5024), .A4(n5025), .Z(n5012) );
  nr03d1 U3034 ( .A1(n5026), .A2(n5027), .A3(n5028), .ZN(n5022) );
  nr04d1 U3035 ( .A1(n5029), .A2(n5030), .A3(n5031), .A4(n5032), .ZN(n5011) );
  nd04d1 U3036 ( .A1(n5033), .A2(n4117), .A3(n4165), .A4(n5036), .ZN(n5029) );
  nr04d1 U3038 ( .A1(n5038), .A2(n5039), .A3(n5040), .A4(n5041), .ZN(n5010) );
  nd12d1 U3040 ( .A1(n5006), .A2(n5045), .ZN(n5009) );
  nr04d1 U3061 ( .A1(n5107), .A2(n5111), .A3(n5112), .A4(n3907), .ZN(n5108) );
  nd04d1 U3119 ( .A1(n5310), .A2(n5304), .A3(n5311), .A4(n4457), .ZN(n5307) );
  nr04d1 U3132 ( .A1(n5352), .A2(n5353), .A3(n4446), .A4(n7152), .ZN(n5351) );
  nr04d1 U3134 ( .A1(n5357), .A2(n4465), .A3(n5358), .A4(n5359), .ZN(n5356) );
  nd04d1 U3137 ( .A1(n5367), .A2(n5368), .A3(n5369), .A4(n3550), .ZN(n5365) );
  nr04d1 U3148 ( .A1(n5401), .A2(n5402), .A3(n5403), .A4(n5404), .ZN(n5400) );
  nr04d1 U3155 ( .A1(n3421), .A2(n6455), .A3(n3331), .A4(n5421), .ZN(n5425) );
  nd04d1 U3160 ( .A1(n3409), .A2(n3410), .A3(n3373), .A4(n5443), .ZN(n5436) );
  nd04d1 U3167 ( .A1(n5463), .A2(n5464), .A3(n3388), .A4(n2807), .ZN(n5460) );
  nd04d1 U3175 ( .A1(n5486), .A2(n5487), .A3(n5488), .A4(n5489), .ZN(n5483) );
  an02d1 U3255 ( .A1(n5638), .A2(n4940), .Z(n5646) );
  nd12d1 U3258 ( .A1(n4942), .A2(n5613), .ZN(n5624) );
  nr03d1 U3259 ( .A1(n5699), .A2(n5700), .A3(n5611), .ZN(n5613) );
  an02d1 U3264 ( .A1(n5590), .A2(n5140), .Z(n5592) );
  an02d1 U3265 ( .A1(n5578), .A2(n4950), .Z(n5590) );
  an03d1 U3270 ( .A1(n4956), .A2(n5706), .A3(n5566), .Z(n5572) );
  nr03d1 U3272 ( .A1(n5708), .A2(n5709), .A3(n5551), .ZN(n5566) );
  an02d1 U3277 ( .A1(n5524), .A2(n5712), .Z(n5536) );
  an02d1 U3280 ( .A1(n4968), .A2(n5511), .Z(n5516) );
  an03d1 U3282 ( .A1(n5380), .A2(n4972), .A3(n5496), .Z(n5508) );
  nr03d1 U3283 ( .A1(n5716), .A2(n12132), .A3(n5493), .ZN(n5496) );
  an02d1 U3288 ( .A1(n5471), .A2(n3266), .Z(n5469) );
  nr03d1 U3289 ( .A1(n4982), .A2(n6670), .A3(n5461), .ZN(n5471) );
  nd04d1 U3290 ( .A1(n3336), .A2(n5721), .A3(n5722), .A4(n5723), .ZN(n5461) );
  nr03d1 U3296 ( .A1(n5726), .A2(n7136), .A3(n5437), .ZN(n5448) );
  nd04d1 U3297 ( .A1(n3337), .A2(n4668), .A3(images_bus[327]), .A4(
        images_bus[324]), .ZN(n5437) );
  nd04d1 U3301 ( .A1(n3480), .A2(n3345), .A3(images_bus[319]), .A4(
        images_bus[316]), .ZN(n5430) );
  an03d1 U3304 ( .A1(n5731), .A2(n5833), .A3(n5408), .Z(n5417) );
  nr04d1 U3305 ( .A1(n3481), .A2(n5733), .A3(n5535), .A4(n6842), .ZN(n5408) );
  nr03d1 U3307 ( .A1(n5636), .A2(n5398), .A3(n5391), .ZN(n5399) );
  nr04d1 U3310 ( .A1(n5373), .A2(n7237), .A3(n6100), .A4(n6173), .ZN(n5375) );
  nd04d1 U3311 ( .A1(n5736), .A2(n4944), .A3(images_bus[285]), .A4(n5413), 
        .ZN(n5373) );
  nr04d1 U3313 ( .A1(n5739), .A2(n5740), .A3(n5741), .A4(n5933), .ZN(n5736) );
  nr04d1 U3314 ( .A1(n5933), .A2(n5742), .A3(n5740), .A4(n5739), .ZN(n5360) );
  nd04d1 U3316 ( .A1(n5743), .A2(n4444), .A3(n4683), .A4(n5349), .ZN(n5739) );
  nr03d1 U3326 ( .A1(n5754), .A2(n5273), .A3(n5755), .ZN(n5285) );
  an02d1 U3332 ( .A1(n5759), .A2(n5226), .Z(n5245) );
  nr04d1 U3333 ( .A1(n3897), .A2(n5218), .A3(n7079), .A4(n5944), .ZN(n5226) );
  nr04d1 U3335 ( .A1(n5760), .A2(n5216), .A3(n6571), .A4(n5186), .ZN(n5222) );
  nd12d1 U3338 ( .A1(n5764), .A2(n5765), .ZN(n5760) );
  nr03d1 U3342 ( .A1(n5169), .A2(n4318), .A3(n5769), .ZN(n5188) );
  nd12d1 U3349 ( .A1(n5148), .A2(n5777), .ZN(n5162) );
  nr03d1 U3356 ( .A1(n5107), .A2(n3982), .A3(n5112), .ZN(n5114) );
  nr03d1 U3360 ( .A1(n5072), .A2(n7093), .A3(n5786), .ZN(n5085) );
  nd04d1 U3364 ( .A1(n5788), .A2(n5789), .A3(n5790), .A4(n5791), .ZN(n5021) );
  nr03d1 U3365 ( .A1(n5792), .A2(n5793), .A3(n4256), .ZN(n5791) );
  nr03d1 U3367 ( .A1(n4238), .A2(n5799), .A3(n5800), .ZN(n5790) );
  nr04d1 U3370 ( .A1(n5807), .A2(n5808), .A3(n5298), .A4(n5809), .ZN(n5804) );
  nr04d1 U3383 ( .A1(n5842), .A2(n5843), .A3(n5844), .A4(n5841), .ZN(n5838) );
  nr04d1 U3395 ( .A1(n5877), .A2(n5878), .A3(n5879), .A4(n5871), .ZN(n5873) );
  nd04d1 U3398 ( .A1(n5889), .A2(n5880), .A3(n5890), .A4(n5891), .ZN(n5887) );
  nd04d1 U3404 ( .A1(n4122), .A2(n5911), .A3(images_bus[107]), .A4(n5912), 
        .ZN(n5907) );
  nr04d1 U3407 ( .A1(n5918), .A2(n5919), .A3(n5908), .A4(n4107), .ZN(n5916) );
  nr04d1 U3425 ( .A1(n5966), .A2(n5967), .A3(n4016), .A4(n4021), .ZN(n5963) );
  nr04d1 U3429 ( .A1(n5973), .A2(n5974), .A3(n5975), .A4(n5976), .ZN(n5972) );
  nd04d1 U3434 ( .A1(images_bus[169]), .A2(n5991), .A3(images_bus[168]), .A4(
        n5992), .ZN(n5990) );
  nr03d1 U3435 ( .A1(n5993), .A2(n5994), .A3(n4422), .ZN(n5992) );
  nd04d1 U3437 ( .A1(n5161), .A2(n5163), .A3(n3938), .A4(n5998), .ZN(n5996) );
  nr03d1 U3441 ( .A1(n6000), .A2(n6259), .A3(n5846), .ZN(n6006) );
  nr04d1 U3450 ( .A1(n6027), .A2(n6028), .A3(n6029), .A4(n6030), .ZN(n6023) );
  nd04d1 U3482 ( .A1(n3576), .A2(n6114), .A3(n5427), .A4(n6116), .ZN(n6112) );
  nd04d1 U3491 ( .A1(n3519), .A2(n5061), .A3(images_bus[277]), .A4(
        images_bus[274]), .ZN(n6144) );
  nd04d1 U3494 ( .A1(n6154), .A2(n3554), .A3(n6156), .A4(n3556), .ZN(n6153) );
  nd04d1 U3496 ( .A1(n3423), .A2(n3473), .A3(n6161), .A4(n3477), .ZN(n6159) );
  nd04d1 U3500 ( .A1(n3430), .A2(n3470), .A3(n6175), .A4(n3469), .ZN(n6171) );
  nd04d1 U3502 ( .A1(n3432), .A2(images_bus[305]), .A3(n6180), .A4(
        images_bus[304]), .ZN(n6178) );
  nd04d1 U3504 ( .A1(n6184), .A2(n3458), .A3(n3459), .A4(n6186), .ZN(n6182) );
  nr03d1 U3513 ( .A1(n6214), .A2(n6215), .A3(n6216), .ZN(n6213) );
  nr04d1 U3539 ( .A1(n6284), .A2(n6285), .A3(n5475), .A4(n6286), .ZN(n6282) );
  nd04d1 U3550 ( .A1(n5486), .A2(n3283), .A3(n6311), .A4(n6312), .ZN(n6309) );
  nr03d1 U3572 ( .A1(n6363), .A2(n6364), .A3(n6365), .ZN(n6359) );
  nd04d1 U3582 ( .A1(n3199), .A2(n6396), .A3(n3195), .A4(n6398), .ZN(n6393) );
  nd04d1 U3585 ( .A1(n3204), .A2(n3195), .A3(n3199), .A4(n6404), .ZN(n6392) );
  nr04d1 U3591 ( .A1(n6421), .A2(n6422), .A3(n3213), .A4(n6424), .ZN(n6420) );
  nr03d1 U3593 ( .A1(n6429), .A2(n6430), .A3(n6431), .ZN(n6427) );
  nd04d1 U3599 ( .A1(n4721), .A2(n6442), .A3(n3041), .A4(n6446), .ZN(n6433) );
  an04d1 U3603 ( .A1(n6454), .A2(n4730), .A3(n6451), .A4(n3052), .Z(n6453) );
  nr03d1 U3619 ( .A1(n2915), .A2(n3017), .A3(n6428), .ZN(n6501) );
  nd12d1 U3640 ( .A1(n6534), .A2(n4936), .ZN(n6535) );
  nr03d1 U3652 ( .A1(n6554), .A2(n4894), .A3(n6483), .ZN(n6494) );
  nr03d1 U3656 ( .A1(n4300), .A2(n4999), .A3(n6471), .ZN(n6477) );
  nd04d1 U3658 ( .A1(n3132), .A2(n5495), .A3(n4411), .A4(n5904), .ZN(n6471) );
  nd04d1 U3664 ( .A1(n3052), .A2(n6451), .A3(n4950), .A4(images_bus[427]), 
        .ZN(n6457) );
  nr03d1 U3665 ( .A1(n4953), .A2(n12140), .A3(n6444), .ZN(n6451) );
  nd04d1 U3670 ( .A1(n6418), .A2(n6579), .A3(n4901), .A4(images_bus[413]), 
        .ZN(n6429) );
  an02d1 U3673 ( .A1(n4901), .A2(n6579), .Z(n6585) );
  an03d1 U3675 ( .A1(n4303), .A2(images_bus[407]), .A3(n6412), .Z(n6418) );
  an03d1 U3676 ( .A1(n5711), .A2(n5035), .A3(n3142), .Z(n6412) );
  nr03d1 U3679 ( .A1(n6591), .A2(n5145), .A3(n6376), .ZN(n6384) );
  nr03d1 U3688 ( .A1(n6597), .A2(n6318), .A3(n6307), .ZN(n6319) );
  an02d1 U3695 ( .A1(n6257), .A2(n5389), .Z(n6269) );
  an02d1 U3697 ( .A1(n3358), .A2(n4983), .Z(n6257) );
  nd12d1 U3701 ( .A1(n6222), .A2(n6602), .ZN(n6233) );
  nr03d1 U3703 ( .A1(n4990), .A2(n4989), .A3(n6208), .ZN(n6227) );
  an02d1 U3705 ( .A1(n6196), .A2(n6603), .Z(n6205) );
  nr04d1 U3707 ( .A1(n6190), .A2(n4526), .A3(n4993), .A4(n6604), .ZN(n6191) );
  nd04d1 U3709 ( .A1(n6605), .A2(n4437), .A3(n6607), .A4(images_bus[298]), 
        .ZN(n6177) );
  nr03d1 U3713 ( .A1(n6608), .A2(n6613), .A3(n6163), .ZN(n6605) );
  nd04d1 U3714 ( .A1(n4485), .A2(images_bus[288]), .A3(n6609), .A4(n6610), 
        .ZN(n6163) );
  nr03d1 U3715 ( .A1(n6100), .A2(n6611), .A3(n6158), .ZN(n6610) );
  nd04d1 U3720 ( .A1(n3520), .A2(n5743), .A3(n6614), .A4(n4444), .ZN(n6135) );
  nr03d1 U3723 ( .A1(n4449), .A2(n6615), .A3(n6616), .ZN(n6131) );
  nr03d1 U3728 ( .A1(n5750), .A2(n5330), .A3(n3692), .ZN(n6114) );
  an03d1 U3738 ( .A1(n6623), .A2(n5271), .A3(n3899), .Z(n6058) );
  an02d1 U3741 ( .A1(n6036), .A2(n6624), .Z(n6044) );
  nr03d1 U3746 ( .A1(n6011), .A2(n6628), .A3(n6626), .ZN(n6026) );
  nd04d1 U3749 ( .A1(n6627), .A2(n3975), .A3(n6629), .A4(n5849), .ZN(n6008) );
  nd04d1 U3753 ( .A1(images_bus[181]), .A2(images_bus[170]), .A3(n5777), .A4(
        n6633), .ZN(n6000) );
  nd04d1 U3755 ( .A1(n6045), .A2(n4711), .A3(n6635), .A4(n6636), .ZN(n5989) );
  nr03d1 U3756 ( .A1(n6938), .A2(n5676), .A3(n5762), .ZN(n6636) );
  nr03d1 U3757 ( .A1(n3974), .A2(n5762), .A3(n6938), .ZN(n5985) );
  nr04d1 U3759 ( .A1(n6637), .A2(n5112), .A3(n3982), .A4(n7244), .ZN(n6635) );
  nr03d1 U3760 ( .A1(n6637), .A2(n3903), .A3(n5112), .ZN(n5977) );
  nd04d1 U3761 ( .A1(n5971), .A2(n4320), .A3(n5441), .A4(images_bus[146]), 
        .ZN(n6637) );
  nd04d1 U3762 ( .A1(n4039), .A2(n6640), .A3(n4034), .A4(n6642), .ZN(n5973) );
  an03d1 U3764 ( .A1(n5969), .A2(n5970), .A3(n6645), .Z(n5971) );
  an03d1 U3765 ( .A1(n5687), .A2(images_bus[140]), .A3(n5962), .Z(n5969) );
  nr03d1 U3766 ( .A1(n3997), .A2(n7173), .A3(n6647), .ZN(n5962) );
  nr03d1 U3770 ( .A1(n6649), .A2(n6650), .A3(n5946), .ZN(n5950) );
  an03d1 U3772 ( .A1(n6652), .A2(images_bus[119]), .A3(n5929), .Z(n5941) );
  an02d1 U3773 ( .A1(n5579), .A2(n5922), .Z(n5929) );
  nr04d1 U3774 ( .A1(n5908), .A2(n4497), .A3(n5918), .A4(n7097), .ZN(n5922) );
  nd04d1 U3780 ( .A1(n5880), .A2(n5890), .A3(n6657), .A4(n5293), .ZN(n5893) );
  nr03d1 U3781 ( .A1(n5871), .A2(n7251), .A3(n4139), .ZN(n5880) );
  nr03d1 U3783 ( .A1(n7042), .A2(n5858), .A3(n5856), .ZN(n5865) );
  nr03d1 U3785 ( .A1(n5844), .A2(n6662), .A3(n5841), .ZN(n5847) );
  nr04d1 U3791 ( .A1(n7574), .A2(n6671), .A3(n6672), .A4(n6673), .ZN(n5795) );
  nd04d1 U3792 ( .A1(n6674), .A2(n4279), .A3(n5314), .A4(n4373), .ZN(n6673) );
  nr03d1 U3793 ( .A1(n6678), .A2(n6679), .A3(n6680), .ZN(n6674) );
  nd04d1 U3800 ( .A1(n5306), .A2(n6697), .A3(n6702), .A4(n6703), .ZN(n6700) );
  nd04d1 U3804 ( .A1(n6715), .A2(n6716), .A3(n6717), .A4(n6718), .ZN(n6712) );
  an04d1 U3805 ( .A1(n6719), .A2(images_bus[48]), .A3(n6720), .A4(n6709), .Z(
        n6718) );
  nr04d1 U3818 ( .A1(n6763), .A2(n6764), .A3(n6765), .A4(n5853), .ZN(n6761) );
  nr03d1 U3820 ( .A1(n6767), .A2(n6768), .A3(n6769), .ZN(n6766) );
  nd04d1 U3832 ( .A1(n5690), .A2(images_bus[105]), .A3(n6798), .A4(n6799), 
        .ZN(n6794) );
  nr04d1 U3852 ( .A1(n6852), .A2(n6853), .A3(n5066), .A4(n4023), .ZN(n6850) );
  nr03d1 U3854 ( .A1(n6858), .A2(n6859), .A3(n6860), .ZN(n6856) );
  nd04d1 U3879 ( .A1(n5170), .A2(n3945), .A3(images_bus[182]), .A4(n6915), 
        .ZN(n6912) );
  nr03d1 U3890 ( .A1(n6941), .A2(n6942), .A3(n4402), .ZN(n6939) );
  nr04d1 U3893 ( .A1(n6949), .A2(n6950), .A3(n5225), .A4(n6951), .ZN(n6947) );
  nr04d1 U3898 ( .A1(n6959), .A2(n6960), .A3(n6250), .A4(n6961), .ZN(n6957) );
  nr04d1 U3900 ( .A1(n6965), .A2(n6966), .A3(n6066), .A4(n3728), .ZN(n6963) );
  nd04d1 U3927 ( .A1(n5345), .A2(n4949), .A3(n7012), .A4(n7021), .ZN(n7018) );
  nr03d1 U3931 ( .A1(n7029), .A2(n6566), .A3(n4450), .ZN(n7033) );
  nd04d1 U3936 ( .A1(n3424), .A2(n7046), .A3(n3476), .A4(n7048), .ZN(n7043) );
  nr03d1 U3953 ( .A1(n7080), .A2(n7086), .A3(n7087), .ZN(n7084) );
  nd04d1 U3957 ( .A1(n7088), .A2(images_bus[309]), .A3(n7095), .A4(n7096), 
        .ZN(n7092) );
  nd04d1 U3959 ( .A1(n5416), .A2(n7101), .A3(n7102), .A4(n7103), .ZN(n7099) );
  nd04d1 U3961 ( .A1(images_bus[317]), .A2(n7107), .A3(n3446), .A4(n7108), 
        .ZN(n7106) );
  nr03d1 U3962 ( .A1(n3444), .A2(n3487), .A3(n7110), .ZN(n7108) );
  nr04d1 U3979 ( .A1(n7149), .A2(n3329), .A3(n7151), .A4(n3274), .ZN(n7148) );
  nd04d1 U3985 ( .A1(n7165), .A2(n3318), .A3(n3323), .A4(n7167), .ZN(n7164) );
  nr03d1 U3987 ( .A1(n7171), .A2(n6306), .A3(n7172), .ZN(n7168) );
  nr04d1 U3994 ( .A1(n7185), .A2(n6597), .A3(n5523), .A4(n7178), .ZN(n7179) );
  nd04d1 U3996 ( .A1(n3293), .A2(n7189), .A3(n7190), .A4(n7191), .ZN(n7186) );
  nd04d1 U3997 ( .A1(n7187), .A2(n5044), .A3(n7192), .A4(n7189), .ZN(n7191) );
  nd04d1 U4001 ( .A1(n7187), .A2(n4305), .A3(n7195), .A4(n5044), .ZN(n7193) );
  nr04d1 U4011 ( .A1(n7213), .A2(n7214), .A3(n7215), .A4(n6365), .ZN(n7212) );
  nd04d1 U4027 ( .A1(n7259), .A2(n3218), .A3(n3037), .A4(n7262), .ZN(n7257) );
  nd04d1 U4054 ( .A1(n7326), .A2(n7327), .A3(n7328), .A4(n7329), .ZN(n7324) );
  nr04d1 U4055 ( .A1(n7330), .A2(n7331), .A3(n7332), .A4(n7333), .ZN(n7329) );
  an02d1 U4065 ( .A1(n7352), .A2(n7353), .Z(n5696) );
  an03d1 U4068 ( .A1(n4824), .A2(n4933), .A3(n7356), .Z(n7328) );
  nd04d1 U4073 ( .A1(n7360), .A2(n5224), .A3(images_bus[448]), .A4(n7302), 
        .ZN(n7314) );
  nd12d1 U4074 ( .A1(n7303), .A2(n2934), .ZN(n7302) );
  an03d1 U4079 ( .A1(n5701), .A2(n4301), .A3(n7285), .Z(n7291) );
  nr03d1 U4080 ( .A1(n6573), .A2(n5702), .A3(n7281), .ZN(n7285) );
  an02d1 U4085 ( .A1(n4730), .A2(n5621), .Z(n4950) );
  nr03d1 U4086 ( .A1(n4953), .A2(n7366), .A3(n3025), .ZN(n7276) );
  nd04d1 U4090 ( .A1(n7252), .A2(n5706), .A3(n4901), .A4(images_bus[415]), 
        .ZN(n7367) );
  nr03d1 U4101 ( .A1(n7375), .A2(n6736), .A3(n7231), .ZN(n7373) );
  an03d1 U4105 ( .A1(n4964), .A2(n5712), .A3(n7226), .Z(n7229) );
  nr03d1 U4106 ( .A1(n5713), .A2(n6366), .A3(n7220), .ZN(n7226) );
  nr03d1 U4109 ( .A1(n4969), .A2(n6595), .A3(n7201), .ZN(n7206) );
  nr03d1 U4111 ( .A1(n5520), .A2(n6597), .A3(n7178), .ZN(n7187) );
  an03d1 U4118 ( .A1(n4656), .A2(n5997), .A3(n7157), .Z(n7170) );
  an03d1 U4119 ( .A1(n5252), .A2(n7146), .A3(n5720), .Z(n7157) );
  nd04d1 U4122 ( .A1(n3353), .A2(n4983), .A3(n7389), .A4(images_bus[344]), 
        .ZN(n7140) );
  nd04d1 U4127 ( .A1(n3354), .A2(n4426), .A3(n5725), .A4(images_bus[337]), 
        .ZN(n7131) );
  nr03d1 U4130 ( .A1(n4989), .A2(n6371), .A3(n7119), .ZN(n7122) );
  nr04d1 U4137 ( .A1(n5416), .A2(n7395), .A3(n7396), .A4(n3488), .ZN(n7394) );
  nr03d1 U4138 ( .A1(n4992), .A2(n7396), .A3(n3488), .ZN(n7392) );
  nr03d1 U4142 ( .A1(n7400), .A2(n7087), .A3(n7080), .ZN(n7088) );
  an02d1 U4148 ( .A1(n7055), .A2(n4677), .Z(n7061) );
  nd04d1 U4151 ( .A1(n7039), .A2(images_bus[287]), .A3(n4944), .A4(n3503), 
        .ZN(n7404) );
  nr04d1 U4153 ( .A1(n7406), .A2(n5740), .A3(n7029), .A4(n7407), .ZN(n7039) );
  nd04d1 U4156 ( .A1(n7026), .A2(n5743), .A3(n5647), .A4(images_bus[267]), 
        .ZN(n7029) );
  nr03d1 U4159 ( .A1(n7411), .A2(n5330), .A3(n3653), .ZN(n7012) );
  nr03d1 U4163 ( .A1(n5296), .A2(n7413), .A3(n6980), .ZN(n6983) );
  an03d1 U4168 ( .A1(n4954), .A2(images_bus[221]), .A3(n6964), .Z(n6962) );
  an02d1 U4169 ( .A1(n6958), .A2(n6623), .Z(n6964) );
  an02d1 U4170 ( .A1(n7416), .A2(n5759), .Z(n6958) );
  nr03d1 U4171 ( .A1(n7417), .A2(n7418), .A3(n5262), .ZN(n6956) );
  nr03d1 U4173 ( .A1(n6944), .A2(n7079), .A3(n7419), .ZN(n7416) );
  nd04d1 U4175 ( .A1(n7420), .A2(n7421), .A3(n7422), .A4(n6940), .ZN(n6944) );
  an03d1 U4177 ( .A1(n5849), .A2(n5435), .A3(n6918), .Z(n6928) );
  nr03d1 U4181 ( .A1(n5774), .A2(n6634), .A3(n6907), .ZN(n6918) );
  nr03d1 U4183 ( .A1(n7429), .A2(n7430), .A3(n7431), .ZN(n6905) );
  nd04d1 U4185 ( .A1(n6881), .A2(n6045), .A3(n4719), .A4(n5683), .ZN(n7431) );
  nr03d1 U4189 ( .A1(n6630), .A2(n5278), .A3(n6876), .ZN(n6881) );
  nr04d1 U4192 ( .A1(n6863), .A2(n5112), .A3(n7434), .A4(n3903), .ZN(n6865) );
  nd04d1 U4193 ( .A1(n6857), .A2(n4320), .A3(n6645), .A4(images_bus[146]), 
        .ZN(n6863) );
  nr03d1 U4194 ( .A1(n5573), .A2(n5952), .A3(n7093), .ZN(n6645) );
  an04d1 U4195 ( .A1(n5970), .A2(n4735), .A3(n6845), .A4(n7435), .Z(n6857) );
  nr03d1 U4196 ( .A1(n7436), .A2(n7173), .A3(n6575), .ZN(n7435) );
  an02d1 U4201 ( .A1(n6836), .A2(n3991), .Z(n6843) );
  nr03d1 U4202 ( .A1(n6650), .A2(n6825), .A3(n4133), .ZN(n6836) );
  nr03d1 U4204 ( .A1(n7034), .A2(n5855), .A3(n6819), .ZN(n6824) );
  an03d1 U4209 ( .A1(n7440), .A2(images_bus[112]), .A3(n6802), .Z(n6808) );
  nr03d1 U4212 ( .A1(n5918), .A2(n7443), .A3(n6796), .ZN(n6802) );
  an03d1 U4214 ( .A1(images_bus[103]), .A2(n6657), .A3(n6784), .Z(n6793) );
  an03d1 U4215 ( .A1(n5890), .A2(n5293), .A3(n6779), .Z(n6784) );
  an04d1 U4217 ( .A1(n4323), .A2(n5852), .A3(n6760), .A4(n7446), .Z(n6772) );
  nr03d1 U4218 ( .A1(n7447), .A2(n6805), .A3(n7042), .ZN(n7446) );
  nd12d1 U4232 ( .A1(n6722), .A2(n7455), .ZN(n6739) );
  nr03d1 U4234 ( .A1(n6589), .A2(n7457), .A3(n6705), .ZN(n6709) );
  nd04d1 U4235 ( .A1(n5306), .A2(n6697), .A3(images_bus[41]), .A4(n6702), .ZN(
        n6705) );
  an03d1 U4240 ( .A1(n4816), .A2(n7466), .A3(n4854), .Z(n7464) );
  nr04d1 U4244 ( .A1(n7479), .A2(n7480), .A3(n7481), .A4(n4334), .ZN(n7475) );
  nr04d1 U4260 ( .A1(n7521), .A2(n7522), .A3(n7523), .A4(n6740), .ZN(n7518) );
  nr04d1 U4265 ( .A1(n7539), .A2(n7540), .A3(n5831), .A4(n7541), .ZN(n7537) );
  nd04d1 U4270 ( .A1(n4207), .A2(n5582), .A3(n7554), .A4(n7555), .ZN(n7550) );
  nd04d1 U4274 ( .A1(n7564), .A2(n7562), .A3(n7565), .A4(n7566), .ZN(n7563) );
  nd04d1 U4275 ( .A1(n6771), .A2(n4065), .A3(n7568), .A4(n4064), .ZN(n7566) );
  nd04d1 U4297 ( .A1(n7614), .A2(n4013), .A3(n6648), .A4(n7616), .ZN(n7613) );
  nd04d1 U4299 ( .A1(n4026), .A2(n7620), .A3(n4052), .A4(n7622), .ZN(n7618) );
  nd04d1 U4305 ( .A1(n7636), .A2(n7637), .A3(n7638), .A4(n7639), .ZN(n7634) );
  nr04d1 U4311 ( .A1(n7651), .A2(n7652), .A3(n7653), .A4(n4424), .ZN(n7649) );
  nd04d1 U4319 ( .A1(n3828), .A2(n7672), .A3(n3835), .A4(n7674), .ZN(n7671) );
  nr03d1 U4320 ( .A1(n6632), .A2(n4390), .A3(n6009), .ZN(n7674) );
  nd04d1 U4324 ( .A1(n3889), .A2(images_bus[201]), .A3(n7685), .A4(
        images_bus[198]), .ZN(n7683) );
  nr03d1 U4328 ( .A1(n7694), .A2(n6571), .A3(n5218), .ZN(n7693) );
  nd04d1 U4332 ( .A1(n3888), .A2(n3859), .A3(n7706), .A4(n7707), .ZN(n7702) );
  nd04d1 U4338 ( .A1(n7718), .A2(n3748), .A3(n3808), .A4(n7720), .ZN(n7717) );
  an03d1 U4342 ( .A1(n3773), .A2(n7725), .A3(n3770), .Z(n7728) );
  an04d1 U4390 ( .A1(n7832), .A2(n7838), .A3(n7839), .A4(n7840), .Z(n7837) );
  nr04d1 U4432 ( .A1(n3124), .A2(n7935), .A3(n5583), .A4(n7936), .ZN(n7933) );
  nr03d1 U4438 ( .A1(n7945), .A2(n7946), .A3(n7366), .ZN(n7944) );
  nr03d1 U4442 ( .A1(n7954), .A2(n3075), .A3(n4406), .ZN(n7953) );
  nr03d1 U4444 ( .A1(n4953), .A2(n7366), .A3(n7945), .ZN(n7932) );
  nd04d1 U4460 ( .A1(n7294), .A2(n2922), .A3(n2946), .A4(n7978), .ZN(n7967) );
  nr04d1 U4461 ( .A1(n7979), .A2(n7313), .A3(n4803), .A4(n5654), .ZN(n7978) );
  nd04d1 U4472 ( .A1(n2877), .A2(n7354), .A3(n2826), .A4(n8004), .ZN(n7995) );
  nr04d1 U4476 ( .A1(n8011), .A2(n8012), .A3(n8013), .A4(n2890), .ZN(n8007) );
  nd12d1 U4481 ( .A1(n8023), .A2(n8024), .ZN(n4911) );
  nd04d1 U4484 ( .A1(n2828), .A2(n2842), .A3(n8029), .A4(n6074), .ZN(n7994) );
  nr03d1 U4485 ( .A1(n8030), .A2(n8031), .A3(n2945), .ZN(n7294) );
  an03d1 U4487 ( .A1(n2922), .A2(n8034), .A3(images_bus[448]), .Z(n7301) );
  nr03d1 U4490 ( .A1(n8040), .A2(n4635), .A3(n2945), .ZN(n8037) );
  nd04d1 U4495 ( .A1(n3015), .A2(n2925), .A3(n2938), .A4(n3009), .ZN(n7309) );
  an02d1 U4504 ( .A1(n8053), .A2(n3109), .Z(n4770) );
  nd12d1 U4506 ( .A1(n7924), .A2(n5729), .ZN(n7945) );
  an03d1 U4517 ( .A1(n5518), .A2(n4961), .A3(n3156), .Z(n7903) );
  nr03d1 U4522 ( .A1(n6591), .A2(n5145), .A3(n7881), .ZN(n7886) );
  nd12d1 U4523 ( .A1(n7876), .A2(n6592), .ZN(n7881) );
  an03d1 U4524 ( .A1(n4967), .A2(n4968), .A3(n5987), .Z(n6592) );
  nd12d1 U4528 ( .A1(n7871), .A2(n4913), .ZN(n8060) );
  an02d1 U4535 ( .A1(n8068), .A2(n4975), .Z(n7864) );
  nr03d1 U4537 ( .A1(n5631), .A2(n5146), .A3(n7855), .ZN(n7860) );
  nd12d1 U4540 ( .A1(n7849), .A2(n5720), .ZN(n7848) );
  an03d1 U4545 ( .A1(n7384), .A2(n3316), .A3(n3277), .Z(n7165) );
  an02d1 U4546 ( .A1(n3339), .A2(n4983), .Z(n7832) );
  nd12d1 U4548 ( .A1(n7830), .A2(n4985), .ZN(n7828) );
  nr03d1 U4551 ( .A1(n4989), .A2(n6371), .A3(n7816), .ZN(n7820) );
  nr03d1 U4554 ( .A1(n4993), .A2(n6604), .A3(n7798), .ZN(n7808) );
  an04d1 U4561 ( .A1(n8075), .A2(n5735), .A3(n6018), .A4(n7777), .Z(n7782) );
  an02d1 U4568 ( .A1(images_bus[264]), .A2(n6134), .Z(n5743) );
  nr04d1 U4570 ( .A1(n7725), .A2(n5750), .A3(n7411), .A4(n5330), .ZN(n7739) );
  nd04d1 U4573 ( .A1(n5655), .A2(images_bus[235]), .A3(n6033), .A4(n8080), 
        .ZN(n7721) );
  nr03d1 U4586 ( .A1(n5186), .A2(n6390), .A3(n5216), .ZN(n7421) );
  nr03d1 U4605 ( .A1(n5062), .A2(n5194), .A3(n7436), .ZN(n5075) );
  nr03d1 U4607 ( .A1(n8100), .A2(n6397), .A3(n5053), .ZN(n5058) );
  nr03d1 U4610 ( .A1(n6650), .A2(n6825), .A3(n7596), .ZN(n7605) );
  nr03d1 U4614 ( .A1(n7442), .A2(n6576), .A3(n7577), .ZN(n7580) );
  nd04d1 U4615 ( .A1(n5690), .A2(n6656), .A3(n4130), .A4(n8102), .ZN(n7577) );
  an03d1 U4616 ( .A1(images_bus[107]), .A2(n5293), .A3(n6657), .Z(n8102) );
  an03d1 U4619 ( .A1(n4117), .A2(n8104), .A3(n8105), .Z(n6771) );
  nr03d1 U4623 ( .A1(n8109), .A2(n7042), .A3(n7559), .ZN(n7562) );
  an03d1 U4633 ( .A1(n5693), .A2(n6665), .A3(n4210), .Z(n7536) );
  nd12d1 U4643 ( .A1(n7512), .A2(n7455), .ZN(n7522) );
  nd04d1 U4647 ( .A1(n6702), .A2(n8119), .A3(images_bus[41]), .A4(n8120), .ZN(
        n7504) );
  an02d1 U4648 ( .A1(n6697), .A2(n4291), .Z(n8120) );
  nd04d1 U4653 ( .A1(n7483), .A2(n8126), .A3(images_bus[28]), .A4(n8127), .ZN(
        n7491) );
  nr03d1 U4654 ( .A1(n7047), .A2(n7481), .A3(n4334), .ZN(n7483) );
  nr04d1 U4656 ( .A1(n8128), .A2(n8129), .A3(n8130), .A4(n7461), .ZN(N26361)
         );
  nr04d1 U4677 ( .A1(n8185), .A2(n7458), .A3(n6690), .A4(n4238), .ZN(n8183) );
  nd04d1 U4683 ( .A1(n8193), .A2(images_bus[45]), .A3(n2793), .A4(n8201), .ZN(
        n8198) );
  nr03d1 U4689 ( .A1(n4255), .A2(n8214), .A3(n8215), .ZN(n8212) );
  an04d1 U4690 ( .A1(n8216), .A2(n4269), .A3(n7455), .A4(n8218), .Z(n8211) );
  an03d1 U4699 ( .A1(n4187), .A2(images_bus[70]), .A3(n5033), .Z(n7529) );
  nd04d1 U4703 ( .A1(n4220), .A2(images_bus[74]), .A3(n8248), .A4(n8249), .ZN(
        n8245) );
  nr04d1 U4707 ( .A1(n4177), .A2(n8258), .A3(n5016), .A4(n8259), .ZN(n8257) );
  nr03d1 U4736 ( .A1(n3996), .A2(n6397), .A3(n8100), .ZN(n8319) );
  nr03d1 U4742 ( .A1(n8331), .A2(n4403), .A3(n8332), .ZN(n8329) );
  nr04d1 U4748 ( .A1(n8348), .A2(n5123), .A3(n5781), .A4(n5117), .ZN(n8347) );
  nr03d1 U4758 ( .A1(n8370), .A2(n8364), .A3(n7081), .ZN(n8368) );
  nr04d1 U4763 ( .A1(n6631), .A2(n8379), .A3(n5184), .A4(n8375), .ZN(n8378) );
  nr03d1 U4774 ( .A1(n8399), .A2(n8400), .A3(n8394), .ZN(n8397) );
  nr03d1 U4776 ( .A1(n8403), .A2(n8404), .A3(n8394), .ZN(n8402) );
  nr04d1 U4807 ( .A1(n8462), .A2(n8463), .A3(n8464), .A4(n8465), .ZN(n8461) );
  nr04d1 U4809 ( .A1(n8467), .A2(n8468), .A3(n4446), .A4(n7754), .ZN(n8466) );
  nr03d1 U4823 ( .A1(n8498), .A2(n8499), .A3(n8492), .ZN(n8494) );
  nd04d1 U4827 ( .A1(n8509), .A2(n7053), .A3(n3468), .A4(n3424), .ZN(n7776) );
  nd12d1 U4836 ( .A1(n8523), .A2(n8524), .ZN(n7074) );
  nr04d1 U4841 ( .A1(n3453), .A2(n8534), .A3(n7085), .A4(n6181), .ZN(n6184) );
  an04d1 U4847 ( .A1(n6194), .A2(n5416), .A3(n3445), .A4(n8539), .Z(n8532) );
  an02d1 U4861 ( .A1(n8564), .A2(n3399), .Z(n5451) );
  nd04d1 U4870 ( .A1(n8580), .A2(n6277), .A3(n8581), .A4(n8582), .ZN(n8576) );
  nd04d1 U4877 ( .A1(n8593), .A2(n6314), .A3(n8594), .A4(n6311), .ZN(n8588) );
  nr03d1 U4884 ( .A1(n8609), .A2(n6997), .A3(n8610), .ZN(n8605) );
  nr04d1 U4889 ( .A1(n8620), .A2(n8621), .A3(n8622), .A4(n8623), .ZN(n8061) );
  nr03d1 U4892 ( .A1(n8629), .A2(n3182), .A3(n3152), .ZN(n8625) );
  nr04d1 U4902 ( .A1(n8653), .A2(n8654), .A3(n8651), .A4(n5562), .ZN(n8652) );
  nr03d1 U4915 ( .A1(n8686), .A2(n7205), .A3(n4955), .ZN(n8685) );
  nr03d1 U4930 ( .A1(n4406), .A2(n3076), .A3(n2796), .ZN(n8710) );
  nr03d1 U4935 ( .A1(n8720), .A2(n3079), .A3(n4408), .ZN(n8719) );
  nd04d1 U4946 ( .A1(n8039), .A2(images_bus[448]), .A3(n8033), .A4(n8038), 
        .ZN(n8743) );
  nd04d1 U4948 ( .A1(n2944), .A2(n3005), .A3(n2948), .A4(n8750), .ZN(n8742) );
  nd04d1 U4956 ( .A1(n7326), .A2(n2983), .A3(n8772), .A4(n8773), .ZN(n8770) );
  nr03d1 U4966 ( .A1(n8796), .A2(n4850), .A3(n2845), .ZN(n7327) );
  nd04d1 U4970 ( .A1(n8803), .A2(n7351), .A3(n8804), .A4(n8805), .ZN(n8799) );
  nr03d1 U4977 ( .A1(n8820), .A2(images_bus[495]), .A3(n8821), .ZN(n8819) );
  nr03d1 U5002 ( .A1(n7375), .A2(n4302), .A3(n8639), .ZN(n8645) );
  an02d1 U5009 ( .A1(n7378), .A2(n8618), .Z(n8619) );
  an03d1 U5011 ( .A1(n4645), .A2(n4968), .A3(images_bus[389]), .Z(n7378) );
  an03d1 U5022 ( .A1(images_bus[376]), .A2(n8608), .A3(n5380), .Z(n8611) );
  nr04d1 U5024 ( .A1(n5716), .A2(n5520), .A3(n7067), .A4(n3259), .ZN(n8604) );
  nr03d1 U5027 ( .A1(n5631), .A2(n4611), .A3(n8589), .ZN(n8593) );
  nd04d1 U5039 ( .A1(images_bus[336]), .A2(n8846), .A3(n4985), .A4(n8847), 
        .ZN(n8568) );
  an02d1 U5040 ( .A1(images_bus[341]), .A2(n6243), .Z(n8847) );
  nr03d1 U5044 ( .A1(n3400), .A2(n8850), .A3(n6237), .ZN(n8564) );
  nr04d1 U5048 ( .A1(n6216), .A2(n7125), .A3(n6226), .A4(images_bus[331]), 
        .ZN(n8851) );
  an03d1 U5051 ( .A1(n7391), .A2(images_bus[326]), .A3(n8542), .Z(n8552) );
  nr03d1 U5052 ( .A1(n6606), .A2(n5254), .A3(n4663), .ZN(n7391) );
  an02d1 U5055 ( .A1(n8535), .A2(n7393), .Z(n8546) );
  nr03d1 U5056 ( .A1(n6098), .A2(n4993), .A3(n4526), .ZN(n7393) );
  an02d1 U5057 ( .A1(n8536), .A2(n5406), .Z(n8535) );
  nr03d1 U5061 ( .A1(n5535), .A2(n8525), .A3(n7400), .ZN(n8529) );
  nr03d1 U5067 ( .A1(n6613), .A2(n5265), .A3(n6608), .ZN(n5735) );
  an02d1 U5068 ( .A1(n8075), .A2(n8503), .Z(n8504) );
  an02d1 U5085 ( .A1(images_bus[248]), .A2(n8856), .Z(n8452) );
  nd04d1 U5086 ( .A1(n8446), .A2(images_bus[247]), .A3(n8857), .A4(n7003), 
        .ZN(n8856) );
  nr03d1 U5089 ( .A1(n7076), .A2(n8441), .A3(n6106), .ZN(n8446) );
  nr03d1 U5090 ( .A1(n8078), .A2(n8858), .A3(n8437), .ZN(n8441) );
  nr03d1 U5094 ( .A1(n7242), .A2(n8428), .A3(n6025), .ZN(n8859) );
  nr03d1 U5101 ( .A1(n4314), .A2(n8863), .A3(n8409), .ZN(n8411) );
  nr03d1 U5107 ( .A1(n5769), .A2(n6631), .A3(n8375), .ZN(n8381) );
  nr03d1 U5109 ( .A1(n7081), .A2(n8364), .A3(n6634), .ZN(n8369) );
  nd12d1 U5114 ( .A1(n6880), .A2(n8867), .ZN(n4424) );
  an04d1 U5115 ( .A1(n5780), .A2(n4725), .A3(images_bus[163]), .A4(n8346), .Z(
        n8350) );
  an02d1 U5123 ( .A1(n5077), .A2(images_bus[139]), .Z(n5970) );
  nr03d1 U5125 ( .A1(n7436), .A2(n6575), .A3(n8318), .ZN(n8324) );
  nd12d1 U5127 ( .A1(n8100), .A2(n8870), .ZN(n6647) );
  nr03d1 U5131 ( .A1(n6649), .A2(n6650), .A3(n8304), .ZN(n8308) );
  nr04d1 U5134 ( .A1(n8873), .A2(n5926), .A3(n7097), .A4(n8296), .ZN(n8300) );
  nr03d1 U5143 ( .A1(n5918), .A2(n7443), .A3(n8878), .ZN(n8283) );
  nd04d1 U5146 ( .A1(n4128), .A2(images_bus[103]), .A3(n6657), .A4(n5293), 
        .ZN(n8879) );
  nr03d1 U5163 ( .A1(n6641), .A2(n5298), .A3(n4751), .ZN(n6666) );
  nr04d1 U5171 ( .A1(n8187), .A2(n6589), .A3(n7457), .A4(n5704), .ZN(n8193) );
  an03d1 U5177 ( .A1(images_bus[28]), .A2(n8127), .A3(n4339), .Z(n8170) );
  nd12d1 U5182 ( .A1(n8888), .A2(n5595), .ZN(n7469) );
  nr04d1 U5184 ( .A1(n8141), .A2(n6355), .A3(n4608), .A4(n6590), .ZN(n8153) );
  nr04d1 U5206 ( .A1(n8930), .A2(n8931), .A3(n8123), .A4(n4346), .ZN(n8927) );
  nd04d1 U5218 ( .A1(n6720), .A2(n8197), .A3(n8955), .A4(n8956), .ZN(n8953) );
  nd04d1 U5221 ( .A1(n4253), .A2(n4259), .A3(n4269), .A4(n8962), .ZN(n8958) );
  nr03d1 U5238 ( .A1(n9003), .A2(n4751), .A3(n8996), .ZN(n8999) );
  nr03d1 U5257 ( .A1(n5882), .A2(n9042), .A3(n4114), .ZN(n9040) );
  nr04d1 U5269 ( .A1(n9066), .A2(n9063), .A3(n9067), .A4(n4135), .ZN(n9065) );
  nd12d1 U5272 ( .A1(n9071), .A2(n9072), .ZN(n5935) );
  nd04d1 U5275 ( .A1(n4098), .A2(n9081), .A3(n4966), .A4(n9082), .ZN(n9079) );
  an02d1 U5292 ( .A1(n5092), .A2(n9115), .Z(n9114) );
  nd12d1 U5326 ( .A1(n5215), .A2(images_bus[204]), .ZN(n9161) );
  nr04d1 U5336 ( .A1(n9184), .A2(n8424), .A3(n6475), .A4(n9185), .ZN(n9183) );
  nr03d1 U5346 ( .A1(n9210), .A2(n9211), .A3(n9212), .ZN(n9209) );
  nr03d1 U5356 ( .A1(n5426), .A2(n9226), .A3(n7017), .ZN(n9230) );
  nr04d1 U5369 ( .A1(n9253), .A2(n6753), .A3(n3541), .A4(n9254), .ZN(n9252) );
  nr03d1 U5396 ( .A1(n9310), .A2(n9309), .A3(n9312), .ZN(n7100) );
  nd04d1 U5398 ( .A1(images_bus[313]), .A2(images_bus[312]), .A3(n9315), .A4(
        n9311), .ZN(n9316) );
  nr04d1 U5409 ( .A1(n3341), .A2(n3409), .A3(n7136), .A4(n5633), .ZN(n9340) );
  an03d1 U5436 ( .A1(n6316), .A2(n6311), .A3(n3283), .Z(n9387) );
  nr04d1 U5458 ( .A1(n9434), .A2(n9435), .A3(n9436), .A4(n9437), .ZN(n9433) );
  nd04d1 U5466 ( .A1(n6579), .A2(n3220), .A3(n7374), .A4(n5806), .ZN(n9446) );
  nr04d1 U5487 ( .A1(n9476), .A2(n9477), .A3(n9478), .A4(n9479), .ZN(n9475) );
  nr04d1 U5501 ( .A1(n9499), .A2(n9500), .A3(n9501), .A4(n8744), .ZN(n9498) );
  an03d1 U5507 ( .A1(n8751), .A2(n5979), .A3(n7315), .Z(n9515) );
  nr03d1 U5530 ( .A1(n8828), .A2(images_bus[492]), .A3(n2910), .ZN(n9560) );
  an03d1 U5542 ( .A1(n9586), .A2(n2868), .A3(n2860), .Z(n9585) );
  nd04d1 U5560 ( .A1(n5380), .A2(images_bus[379]), .A3(images_bus[376]), .A4(
        n9405), .ZN(n9605) );
  an03d1 U5563 ( .A1(images_bus[368]), .A2(n9392), .A3(n4975), .Z(n9397) );
  nd12d1 U5566 ( .A1(n9391), .A2(n8070), .ZN(n9392) );
  nd04d1 U5569 ( .A1(n7382), .A2(images_bus[363]), .A3(images_bus[360]), .A4(
        n9385), .ZN(n9608) );
  an02d1 U5574 ( .A1(images_bus[348]), .A2(n9609), .Z(n9371) );
  nd04d1 U5575 ( .A1(n7388), .A2(images_bus[347]), .A3(images_bus[344]), .A4(
        n3342), .ZN(n9609) );
  an03d1 U5588 ( .A1(n9610), .A2(n3409), .A3(n3405), .Z(n7818) );
  nd04d1 U5590 ( .A1(n5634), .A2(images_bus[331]), .A3(images_bus[328]), .A4(
        n9341), .ZN(n9611) );
  an02d1 U5600 ( .A1(n9320), .A2(n3345), .Z(n9321) );
  an02d1 U5614 ( .A1(n9283), .A2(n4677), .Z(n9287) );
  an02d1 U5621 ( .A1(n9267), .A2(n3503), .Z(n9272) );
  nd12d1 U5628 ( .A1(n9620), .A2(images_bus[272]), .ZN(n5740) );
  an03d1 U5629 ( .A1(images_bus[264]), .A2(n9244), .A3(n5647), .Z(n9251) );
  an02d1 U5633 ( .A1(n5345), .A2(images_bus[255]), .Z(n6617) );
  nr04d1 U5635 ( .A1(n7411), .A2(n7017), .A3(n4948), .A4(n9226), .ZN(n9622) );
  nr03d1 U5642 ( .A1(n9201), .A2(n12118), .A3(n7413), .ZN(n9211) );
  nr03d1 U5648 ( .A1(n6025), .A2(n9197), .A3(n3719), .ZN(n9201) );
  nr03d1 U5657 ( .A1(n7079), .A2(n9169), .A3(n5234), .ZN(n9173) );
  nr03d1 U5658 ( .A1(n5218), .A2(n5944), .A3(n9163), .ZN(n9169) );
  nd04d1 U5660 ( .A1(n8401), .A2(images_bus[203]), .A3(images_bus[200]), .A4(
        n9628), .ZN(n9627) );
  nd12d1 U5668 ( .A1(n9145), .A2(n5767), .ZN(n9151) );
  nd12d1 U5671 ( .A1(n9137), .A2(n8865), .ZN(n9143) );
  nd04d1 U5673 ( .A1(n5567), .A2(images_bus[176]), .A3(images_bus[179]), .A4(
        n9136), .ZN(n9630) );
  an02d1 U5676 ( .A1(n9132), .A2(n3932), .Z(n7654) );
  an03d1 U5677 ( .A1(n3927), .A2(n6902), .A3(n3928), .Z(n9132) );
  an02d1 U5689 ( .A1(n9115), .A2(n5783), .Z(n9113) );
  an02d1 U5692 ( .A1(images_bus[140]), .A2(n9637), .Z(n9102) );
  nd04d1 U5693 ( .A1(n5687), .A2(images_bus[139]), .A3(images_bus[136]), .A4(
        n9099), .ZN(n9637) );
  nd04d1 U5711 ( .A1(n5690), .A2(images_bus[107]), .A3(images_bus[104]), .A4(
        n9048), .ZN(n9641) );
  nd04d1 U5716 ( .A1(images_bus[91]), .A2(n5458), .A3(images_bus[88]), .A4(
        n9027), .ZN(n9642) );
  nr04d1 U5750 ( .A1(n8907), .A2(n5964), .A3(n6355), .A4(n4608), .ZN(n8920) );
  nd12d1 U5752 ( .A1(n8139), .A2(images_bus[11]), .ZN(n8141) );
  nr03d1 U5781 ( .A1(n9696), .A2(n9697), .A3(n4231), .ZN(n7498) );
  nd04d1 U5794 ( .A1(n4268), .A2(n4262), .A3(n9726), .A4(n9727), .ZN(n9722) );
  an03d1 U5802 ( .A1(n4186), .A2(n4183), .A3(n5033), .Z(n6744) );
  nr04d1 U5816 ( .A1(images_bus[94]), .A2(n9776), .A3(n9777), .A4(n5027), .ZN(
        n9774) );
  nd04d1 U5841 ( .A1(n4391), .A2(n4007), .A3(images_bus[132]), .A4(n9822), 
        .ZN(n9818) );
  nr04d1 U5862 ( .A1(n9865), .A2(n3926), .A3(n6893), .A4(n6889), .ZN(n9864) );
  nd04d1 U5895 ( .A1(n4412), .A2(n3861), .A3(n3870), .A4(n9926), .ZN(n9920) );
  nd12d1 U5920 ( .A1(n5339), .A2(n5338), .ZN(n4410) );
  nr04d1 U5921 ( .A1(n9968), .A2(n9969), .A3(n4948), .A4(n3587), .ZN(n9966) );
  nr04d1 U5958 ( .A1(n10035), .A2(n7090), .A3(n8534), .A4(n9310), .ZN(n10034)
         );
  nd04d1 U6008 ( .A1(n6331), .A2(n3301), .A3(n10108), .A4(n10109), .ZN(n10107)
         );
  nr03d1 U6011 ( .A1(n6593), .A2(n10114), .A3(n6353), .ZN(n10113) );
  nd04d1 U6035 ( .A1(n7259), .A2(n3218), .A3(n3229), .A4(n10159), .ZN(n10158)
         );
  nr03d1 U6038 ( .A1(n8679), .A2(n10167), .A3(n3038), .ZN(n10166) );
  nr04d1 U6076 ( .A1(N14866), .A2(n10240), .A3(n2999), .A4(n2917), .ZN(n10239)
         );
  nd04d1 U6082 ( .A1(n2966), .A2(n2964), .A3(n2993), .A4(n10255), .ZN(n10250)
         );
  nr03d1 U6095 ( .A1(n7335), .A2(n8796), .A3(n7337), .ZN(n9551) );
  nd04d1 U6106 ( .A1(n2877), .A2(n2876), .A3(n2871), .A4(n10309), .ZN(n10306)
         );
  nr03d1 U6125 ( .A1(n6979), .A2(n2896), .A3(n5320), .ZN(n9583) );
  an02d1 U6128 ( .A1(images_bus[502]), .A2(n10323), .Z(n10332) );
  nr03d1 U6132 ( .A1(n10325), .A2(n2891), .A3(n10348), .ZN(n8818) );
  nd12d1 U6133 ( .A1(n10349), .A2(n2878), .ZN(n10325) );
  an02d1 U6149 ( .A1(n10276), .A2(images_bus[479]), .Z(n10277) );
  nd12d1 U6156 ( .A1(n10268), .A2(images_bus[471]), .ZN(n10273) );
  nd04d1 U6160 ( .A1(n2971), .A2(n2979), .A3(n8781), .A4(n6655), .ZN(n10265)
         );
  nr03d1 U6171 ( .A1(n6555), .A2(n10248), .A3(n4397), .ZN(n10245) );
  nr03d1 U6172 ( .A1(n2918), .A2(n12129), .A3(n5126), .ZN(n10248) );
  nr04d1 U6174 ( .A1(n2966), .A2(n10368), .A3(n5484), .A4(n10369), .ZN(n10365)
         );
  nd12d1 U6188 ( .A1(n8740), .A2(n8738), .ZN(n9497) );
  an02d1 U6192 ( .A1(n10220), .A2(images_bus[447]), .Z(n10217) );
  nd12d1 U6196 ( .A1(n10212), .A2(images_bus[443]), .ZN(n10211) );
  nr03d1 U6214 ( .A1(n10384), .A2(n8695), .A3(n4744), .ZN(n10189) );
  an02d1 U6219 ( .A1(n10179), .A2(images_bus[423]), .Z(n10184) );
  nr03d1 U6226 ( .A1(n6160), .A2(n10169), .A3(n6084), .ZN(n10167) );
  an03d1 U6233 ( .A1(n10387), .A2(n6437), .A3(images_bus[413]), .Z(n10169) );
  an02d1 U6242 ( .A1(n10131), .A2(images_bus[395]), .Z(n10137) );
  nr03d1 U6257 ( .A1(n10392), .A2(n12124), .A3(n5242), .ZN(n10390) );
  nr03d1 U6259 ( .A1(n6162), .A2(n10115), .A3(n6089), .ZN(n10118) );
  an03d1 U6262 ( .A1(images_bus[380]), .A2(n10112), .A3(images_bus[381]), .Z(
        n10115) );
  an02d1 U6265 ( .A1(n6295), .A2(n5480), .Z(n6299) );
  an02d1 U6285 ( .A1(n10035), .A2(images_bus[311]), .Z(n10038) );
  an02d1 U6290 ( .A1(n10030), .A2(images_bus[303]), .Z(n10029) );
  nr03d1 U6294 ( .A1(n6842), .A2(n10022), .A3(n5164), .ZN(n10025) );
  nr03d1 U6295 ( .A1(n7150), .A2(n10018), .A3(n5636), .ZN(n10022) );
  nr03d1 U6296 ( .A1(n10016), .A2(n12153), .A3(n6007), .ZN(n10018) );
  nr03d1 U6298 ( .A1(n6613), .A2(n10012), .A3(n4675), .ZN(n10016) );
  an02d1 U6299 ( .A1(n10014), .A2(images_bus[291]), .Z(n10012) );
  nr03d1 U6304 ( .A1(n6173), .A2(n3484), .A3(n6100), .ZN(n10007) );
  nd12d1 U6315 ( .A1(n9987), .A2(images_bus[267]), .ZN(n9986) );
  nd04d1 U6318 ( .A1(n3561), .A2(n5002), .A3(n3562), .A4(n10400), .ZN(n7037)
         );
  an02d1 U6319 ( .A1(n3525), .A2(n10402), .Z(n7027) );
  an02d1 U6331 ( .A1(n9950), .A2(images_bus[239]), .Z(n9951) );
  an02d1 U6344 ( .A1(n9930), .A2(images_bus[219]), .Z(n9928) );
  nr03d1 U6367 ( .A1(n6259), .A2(n9883), .A3(n5846), .ZN(n9884) );
  nr03d1 U6382 ( .A1(n6185), .A2(n9853), .A3(n6123), .ZN(n9850) );
  an02d1 U6396 ( .A1(n9832), .A2(images_bus[143]), .Z(n9830) );
  nd12d1 U6400 ( .A1(n9827), .A2(images_bus[135]), .ZN(n9826) );
  nr03d1 U6406 ( .A1(n6189), .A2(n9815), .A3(n6133), .ZN(n9816) );
  an02d1 U6408 ( .A1(images_bus[122]), .A2(n10417), .Z(n9812) );
  nr03d1 U6420 ( .A1(n5041), .A2(n5015), .A3(n5006), .ZN(n8307) );
  an02d1 U6430 ( .A1(n10421), .A2(n6699), .Z(n9767) );
  nr03d1 U6438 ( .A1(n6882), .A2(n9752), .A3(n5204), .ZN(n9753) );
  an02d1 U6439 ( .A1(n5697), .A2(n9744), .Z(n9752) );
  an02d1 U6452 ( .A1(n10423), .A2(n9008), .Z(n5033) );
  an02d1 U6454 ( .A1(n9715), .A2(images_bus[51]), .Z(n9719) );
  nr03d1 U6457 ( .A1(n6348), .A2(n9712), .A3(n5959), .ZN(n9713) );
  an03d1 U6458 ( .A1(images_bus[44]), .A2(n9708), .A3(images_bus[45]), .Z(
        n9712) );
  an02d1 U6467 ( .A1(n5788), .A2(n10426), .Z(n7500) );
  nr03d1 U6485 ( .A1(n9661), .A2(n10430), .A3(n7588), .ZN(n7466) );
  nd04d1 U6488 ( .A1(n9651), .A2(n5794), .A3(n10433), .A4(images_bus[2]), .ZN(
        n10432) );
  nr03d1 U6507 ( .A1(n9691), .A2(n10471), .A3(n10472), .ZN(n10470) );
  an03d1 U6517 ( .A1(n8197), .A2(n4512), .A3(N8510), .Z(n8950) );
  nd04d1 U6528 ( .A1(n4146), .A2(n4188), .A3(n5779), .A4(n10519), .ZN(n10516)
         );
  nd04d1 U6533 ( .A1(n4150), .A2(n5821), .A3(n9008), .A4(n10530), .ZN(n10528)
         );
  an02d1 U6545 ( .A1(n10542), .A2(n5581), .Z(n5842) );
  an02d1 U6552 ( .A1(n8104), .A2(n4167), .Z(n5872) );
  nr03d1 U6599 ( .A1(n9100), .A2(n5967), .A3(n8323), .ZN(n7620) );
  nr03d1 U6648 ( .A1(n3959), .A2(n3906), .A3(n10661), .ZN(n10659) );
  nd04d1 U6672 ( .A1(n3850), .A2(n10683), .A3(n10684), .A4(n3843), .ZN(n10682)
         );
  nr04d1 U6676 ( .A1(n10692), .A2(n5239), .A3(n8863), .A4(n9919), .ZN(n10691)
         );
  an02d1 U6678 ( .A1(n3854), .A2(n5232), .Z(n8413) );
  an02d1 U6696 ( .A1(n3770), .A2(n8440), .Z(n4420) );
  nr04d1 U6699 ( .A1(n10727), .A2(n6619), .A3(n10728), .A4(n6094), .ZN(n10725)
         );
  an03d1 U6715 ( .A1(images_bus[258]), .A2(n10761), .A3(n8464), .Z(n10760) );
  nd04d1 U6716 ( .A1(n3570), .A2(n10762), .A3(n8468), .A4(n10763), .ZN(n10757)
         );
  nr03d1 U6725 ( .A1(n9254), .A2(n10776), .A3(n5358), .ZN(n10775) );
  nd04d1 U6735 ( .A1(n10794), .A2(n5379), .A3(n10795), .A4(n10796), .ZN(n10793) );
  nr03d1 U6736 ( .A1(n10003), .A2(n5371), .A3(n3555), .ZN(n10796) );
  nd04d1 U6737 ( .A1(n3549), .A2(n3553), .A3(n10795), .A4(n10799), .ZN(n10792)
         );
  nr03d1 U6740 ( .A1(n9273), .A2(n10804), .A3(n9276), .ZN(n10803) );
  nd04d1 U6744 ( .A1(n3473), .A2(n3474), .A3(n6169), .A4(n10811), .ZN(n10810)
         );
  nd04d1 U6749 ( .A1(n3471), .A2(n3469), .A3(n10020), .A4(n10816), .ZN(n10815)
         );
  nr03d1 U6751 ( .A1(n5393), .A2(n10819), .A3(n3431), .ZN(n10818) );
  nd04d1 U6753 ( .A1(n3465), .A2(n10823), .A3(n10824), .A4(n9294), .ZN(n10822)
         );
  nr04d1 U6788 ( .A1(n10868), .A2(n10863), .A3(n10869), .A4(n9336), .ZN(n10867) );
  nr03d1 U6791 ( .A1(n7125), .A2(n10873), .A3(n3406), .ZN(n10872) );
  nr03d1 U6794 ( .A1(n10077), .A2(n10881), .A3(n10882), .ZN(n10880) );
  nr03d1 U6811 ( .A1(n10905), .A2(n3391), .A3(n6275), .ZN(n10904) );
  nr04d1 U6815 ( .A1(n10908), .A2(n3328), .A3(n10910), .A4(n5474), .ZN(n10902)
         );
  nr04d1 U6821 ( .A1(n10923), .A2(n3278), .A3(n7386), .A4(n7385), .ZN(n10922)
         );
  an04d1 U6839 ( .A1(n6353), .A2(n10946), .A3(n6342), .A4(n3305), .Z(n10945)
         );
  nd04d1 U6848 ( .A1(n10958), .A2(images_bus[380]), .A3(n6593), .A4(n10946), 
        .ZN(n10957) );
  nr03d1 U6858 ( .A1(n7225), .A2(n10979), .A3(n6380), .ZN(n10978) );
  nr04d1 U6860 ( .A1(n7889), .A2(n10983), .A3(n10984), .A4(n7884), .ZN(n10982)
         );
  nr04d1 U6873 ( .A1(n11008), .A2(n11009), .A3(n11010), .A4(n7915), .ZN(n11007) );
  nd04d1 U6907 ( .A1(n3111), .A2(n3090), .A3(n11055), .A4(n6486), .ZN(n11054)
         );
  nd04d1 U6910 ( .A1(n3095), .A2(n3106), .A3(n11061), .A4(n11062), .ZN(n11060)
         );
  nd04d1 U6924 ( .A1(n2937), .A2(n2940), .A3(n3011), .A4(n11079), .ZN(n11074)
         );
  an02d1 U6938 ( .A1(images_bus[460]), .A2(n7336), .Z(n10247) );
  nd04d1 U6939 ( .A1(n2989), .A2(n2992), .A3(n2967), .A4(n11095), .ZN(n11090)
         );
  nd12d1 U6948 ( .A1(n9526), .A2(n2973), .ZN(n9528) );
  nd12d1 U6949 ( .A1(n10362), .A2(n10257), .ZN(n9526) );
  nr03d1 U6957 ( .A1(n2842), .A2(n12161), .A3(n11123), .ZN(n11122) );
  nd04d1 U6971 ( .A1(n2872), .A2(n2879), .A3(n2815), .A4(n10350), .ZN(n11147)
         );
  an02d1 U6985 ( .A1(n2888), .A2(n11175), .Z(n9577) );
  nr03d1 U6988 ( .A1(n11174), .A2(N15586), .A3(n11180), .ZN(n11179) );
  an02d1 U6990 ( .A1(images_bus[507]), .A2(n11174), .Z(n11176) );
  nd12d1 U6999 ( .A1(n10333), .A2(n10329), .ZN(n9581) );
  nr03d1 U7018 ( .A1(n11189), .A2(n2868), .A3(n11136), .ZN(n8005) );
  an02d1 U7026 ( .A1(n11193), .A2(n9554), .Z(n9591) );
  nd12d1 U7067 ( .A1(n11087), .A2(n8047), .ZN(n10370) );
  nr04d1 U7073 ( .A1(n9502), .A2(n6894), .A3(n9501), .A4(n8744), .ZN(n11207)
         );
  nr04d1 U7088 ( .A1(n6480), .A2(n6478), .A3(n11056), .A4(n11053), .ZN(n8716)
         );
  an02d1 U7105 ( .A1(images_bus[422]), .A2(n11023), .Z(n11021) );
  an03d1 U7126 ( .A1(n3223), .A2(n6588), .A3(images_bus[408]), .Z(n11218) );
  an02d1 U7175 ( .A1(n8839), .A2(n3301), .Z(n5505) );
  nd04d1 U7182 ( .A1(n6314), .A2(n3281), .A3(n3269), .A4(n11229), .ZN(n10926)
         );
  an02d1 U7216 ( .A1(images_bus[324]), .A2(n10864), .Z(n11236) );
  an02d1 U7219 ( .A1(images_bus[318]), .A2(n10851), .Z(n11237) );
  an02d1 U7260 ( .A1(n4946), .A2(n10790), .Z(n10801) );
  nr03d1 U7275 ( .A1(n6615), .A2(n11243), .A3(n9998), .ZN(n11246) );
  an02d1 U7291 ( .A1(n3526), .A2(n11250), .Z(n10403) );
  nd04d1 U7292 ( .A1(n7751), .A2(n11251), .A3(n11252), .A4(n10761), .ZN(n10751) );
  an02d1 U7308 ( .A1(n3800), .A2(n10407), .Z(n9624) );
  an02d1 U7311 ( .A1(images_bus[240]), .A2(n10724), .Z(n10731) );
  nd12d1 U7319 ( .A1(n9207), .A2(n3761), .ZN(n4407) );
  nd12d1 U7347 ( .A1(n5227), .A2(n5219), .ZN(n6950) );
  an02d1 U7419 ( .A1(n6821), .A2(n4085), .Z(n5036) );
  an02d1 U7429 ( .A1(images_bus[104]), .A2(n10561), .Z(n10565) );
  nr03d1 U7447 ( .A1(n11283), .A2(images_bus[91]), .A3(n5866), .ZN(n8881) );
  nd12d1 U7466 ( .A1(n6765), .A2(n10542), .ZN(n5848) );
  an02d1 U7503 ( .A1(images_bus[30]), .A2(n10469), .Z(n10476) );
  an02d1 U7510 ( .A1(images_bus[23]), .A2(n11296), .Z(n10462) );
  nr03d1 U7529 ( .A1(n8129), .A2(n8137), .A3(n11300), .ZN(n7463) );
  nr03d1 U7531 ( .A1(n7574), .A2(n5785), .A3(n5008), .ZN(n9651) );
  nd04d1 U7536 ( .A1(N8008), .A2(n5794), .A3(n11304), .A4(n11305), .ZN(n11303)
         );
  an02d1 U7545 ( .A1(N8074), .A2(n4844), .Z(n8131) );
  an02d1 U7548 ( .A1(N8054), .A2(n4847), .Z(n8900) );
  nr03d1 U7566 ( .A1(n9670), .A2(images_bus[19]), .A3(n8909), .ZN(n7471) );
  nr04d1 U7595 ( .A1(n11334), .A2(n11335), .A3(n8168), .A4(n7494), .ZN(n11332)
         );
  nr03d1 U7596 ( .A1(n8171), .A2(n11336), .A3(n9687), .ZN(n7494) );
  nd12d1 U7603 ( .A1(n10472), .A2(N8330), .ZN(n8178) );
  nr03d1 U7606 ( .A1(n11340), .A2(n4277), .A3(n6668), .ZN(n11337) );
  an03d1 U7623 ( .A1(n4275), .A2(images_bus[39]), .A3(N8445), .Z(n10489) );
  an02d1 U7624 ( .A1(N8432), .A2(n4275), .Z(n10480) );
  nr04d1 U7633 ( .A1(n11360), .A2(n11361), .A3(n7105), .A4(n7513), .ZN(n11359)
         );
  nd12d1 U7634 ( .A1(n6724), .A2(n6720), .ZN(n7513) );
  an02d1 U7652 ( .A1(N8627), .A2(n4260), .Z(n8967) );
  an03d1 U7653 ( .A1(images_bus[54]), .A2(n4260), .A3(N8640), .Z(n11372) );
  an02d1 U7654 ( .A1(N8653), .A2(n11375), .Z(n9726) );
  nd12d1 U7655 ( .A1(n10508), .A2(n7511), .ZN(n9718) );
  nd04d1 U7658 ( .A1(n4270), .A2(N8575), .A3(n6720), .A4(images_bus[49]), .ZN(
        n8208) );
  nd12d1 U7661 ( .A1(n8964), .A2(n4259), .ZN(n10508) );
  an03d1 U7666 ( .A1(n4269), .A2(n7455), .A3(N8614), .Z(n8216) );
  nd04d1 U7673 ( .A1(n4328), .A2(n11380), .A3(n4228), .A4(n11382), .ZN(n11376)
         );
  an02d1 U7678 ( .A1(n8983), .A2(n8986), .Z(n6734) );
  nd12d1 U7685 ( .A1(n8986), .A2(n8983), .ZN(n8116) );
  an03d1 U7686 ( .A1(n9731), .A2(images_bus[59]), .A3(N8705), .Z(n8983) );
  an02d1 U7687 ( .A1(N8692), .A2(n4266), .Z(n9731) );
  an02d1 U7689 ( .A1(n8991), .A2(n4201), .Z(n8228) );
  an02d1 U7690 ( .A1(n4224), .A2(n9733), .Z(n8991) );
  an03d1 U7691 ( .A1(n8988), .A2(n8884), .A3(N8744), .Z(n9733) );
  nd12d1 U7699 ( .A1(n5809), .A2(N8812), .ZN(n5812) );
  an02d1 U7701 ( .A1(N8826), .A2(n11392), .Z(n10423) );
  an03d1 U7717 ( .A1(n4181), .A2(images_bus[75]), .A3(N8924), .Z(n5829) );
  nd12d1 U7727 ( .A1(n6764), .A2(N9008), .ZN(n6765) );
  an03d1 U7756 ( .A1(n11430), .A2(images_bus[94]), .A3(N9190), .Z(n9032) );
  nd12d1 U7774 ( .A1(n5899), .A2(N9302), .ZN(n5897) );
  an02d1 U7780 ( .A1(N9344), .A2(n6790), .Z(n5909) );
  nr04d1 U7781 ( .A1(n4074), .A2(n11447), .A3(n5689), .A4(n11448), .ZN(n11445)
         );
  an02d1 U7785 ( .A1(N9372), .A2(n5911), .Z(n5914) );
  nd04d1 U7799 ( .A1(n11454), .A2(n6815), .A3(n5579), .A4(n11460), .ZN(n11459)
         );
  an02d1 U7809 ( .A1(N9526), .A2(n4099), .Z(n9076) );
  nr03d1 U7810 ( .A1(n11464), .A2(n7034), .A3(n11462), .ZN(n11463) );
  nd12d1 U7842 ( .A1(n6853), .A2(n9098), .ZN(n8320) );
  an02d1 U7847 ( .A1(N9816), .A2(n4024), .Z(n10603) );
  nd12d1 U7849 ( .A1(n9100), .A2(n4022), .ZN(n5074) );
  an02d1 U7859 ( .A1(N9891), .A2(n4052), .Z(n11275) );
  nr03d1 U7864 ( .A1(n11503), .A2(n5573), .A3(n7093), .ZN(n11502) );
  an03d1 U7871 ( .A1(n4050), .A2(n4319), .A3(N9966), .Z(n7635) );
  an02d1 U7884 ( .A1(N10071), .A2(n4045), .Z(n6640) );
  an02d1 U7889 ( .A1(n4043), .A2(n9848), .Z(n7647) );
  an03d1 U7890 ( .A1(n4044), .A2(images_bus[157]), .A3(N10101), .Z(n9848) );
  nd04d1 U7933 ( .A1(n11536), .A2(n5192), .A3(images_bus[173]), .A4(n11537), 
        .ZN(n11535) );
  an03d1 U7935 ( .A1(n6902), .A2(images_bus[173]), .A3(N10341), .Z(n5157) );
  nd04d1 U7938 ( .A1(n11536), .A2(n5777), .A3(n11539), .A4(n7659), .ZN(n11538)
         );
  an02d1 U8008 ( .A1(N10791), .A2(n9167), .Z(n10683) );
  an02d1 U8030 ( .A1(n3865), .A2(n5257), .Z(n7708) );
  an02d1 U8032 ( .A1(n6055), .A2(n3862), .Z(n6053) );
  nd12d1 U8038 ( .A1(n5264), .A2(n5257), .ZN(n10700) );
  an02d1 U8039 ( .A1(N11031), .A2(n3864), .Z(n5257) );
  an02d1 U8041 ( .A1(n3858), .A2(n11583), .Z(n6055) );
  nd04d1 U8043 ( .A1(n8417), .A2(N11001), .A3(n3861), .A4(images_bus[217]), 
        .ZN(n5262) );
  an02d1 U8044 ( .A1(N10986), .A2(n3861), .Z(n8417) );
  an02d1 U8062 ( .A1(N11166), .A2(n9199), .Z(n6073) );
  an04d1 U8113 ( .A1(n8857), .A2(n7003), .A3(n7743), .A4(n3783), .Z(n6110) );
  nd12d1 U8135 ( .A1(n7015), .A2(N11526), .ZN(n9235) );
  an02d1 U8138 ( .A1(n8453), .A2(images_bus[251]), .Z(n5338) );
  an02d1 U8142 ( .A1(N11571), .A2(n3571), .Z(n11250) );
  an02d1 U8144 ( .A1(n11251), .A2(n5746), .Z(n4435) );
  nd12d1 U8146 ( .A1(n11252), .A2(n11251), .ZN(n4443) );
  an02d1 U8147 ( .A1(N11586), .A2(n3527), .Z(n11251) );
  nd12d1 U8153 ( .A1(n10764), .A2(n11637), .ZN(n9239) );
  nd04d1 U8154 ( .A1(N11650), .A2(n10402), .A3(images_bus[259]), .A4(
        images_bus[260]), .ZN(n10764) );
  nd04d1 U8191 ( .A1(n11656), .A2(n4485), .A3(n11659), .A4(n11660), .ZN(n11658) );
  nd12d1 U8210 ( .A1(n10828), .A2(n11668), .ZN(n7078) );
  an02d1 U8219 ( .A1(n11677), .A2(n7789), .Z(n11676) );
  nr03d1 U8236 ( .A1(n8534), .A2(n3452), .A3(n9310), .ZN(n7792) );
  nd12d1 U8246 ( .A1(n9304), .A2(N12434), .ZN(n9310) );
  nd12d1 U8253 ( .A1(n9315), .A2(n6194), .ZN(n4517) );
  nr04d1 U8257 ( .A1(n11692), .A2(n4535), .A3(n4536), .A4(n11693), .ZN(n11691)
         );
  nd12d1 U8281 ( .A1(n10067), .A2(n3408), .ZN(n11708) );
  nd04d1 U8291 ( .A1(n4986), .A2(n4987), .A3(n11711), .A4(n11713), .ZN(n11712)
         );
  an02d1 U8293 ( .A1(n3377), .A2(n11716), .Z(n4563) );
  nd04d1 U8303 ( .A1(n6263), .A2(n3395), .A3(n11720), .A4(n5397), .ZN(n11725)
         );
  an02d1 U8306 ( .A1(n3396), .A2(n11723), .Z(n11720) );
  nd12d1 U8310 ( .A1(n5455), .A2(N12946), .ZN(n6258) );
  nr04d1 U8316 ( .A1(n4570), .A2(n11727), .A3(n3384), .A4(n11719), .ZN(n11717)
         );
  nr03d1 U8319 ( .A1(n3387), .A2(n5721), .A3(n11721), .ZN(n11728) );
  nd12d1 U8348 ( .A1(n9379), .A2(N13202), .ZN(n6301) );
  an02d1 U8371 ( .A1(n10935), .A2(n5523), .Z(n4620) );
  nd12d1 U8377 ( .A1(n10106), .A2(n7189), .ZN(n11765) );
  an03d1 U8381 ( .A1(n3312), .A2(n5504), .A3(n7189), .Z(n8067) );
  nd12d1 U8384 ( .A1(n8066), .A2(n5719), .ZN(n4630) );
  an02d1 U8388 ( .A1(n4972), .A2(n7198), .Z(n4627) );
  nr03d1 U8410 ( .A1(n8842), .A2(n11779), .A3(n10120), .ZN(n8063) );
  an02d1 U8443 ( .A1(n3243), .A2(n8626), .Z(n11794) );
  nd04d1 U8463 ( .A1(n11219), .A2(n3239), .A3(n6416), .A4(n4302), .ZN(n11810)
         );
  an02d1 U8473 ( .A1(N13938), .A2(n11220), .Z(n11219) );
  nr04d1 U8477 ( .A1(n6588), .A2(n8057), .A3(n3220), .A4(images_bus[409]), 
        .ZN(n11812) );
  nr03d1 U8484 ( .A1(n6430), .A2(images_bus[413]), .A3(n6431), .ZN(n11818) );
  nr03d1 U8504 ( .A1(n3051), .A2(images_bus[419]), .A3(n6577), .ZN(n4718) );
  nd04d1 U8511 ( .A1(n3127), .A2(n3054), .A3(n11828), .A4(n5980), .ZN(n11827)
         );
  nr03d1 U8516 ( .A1(n7935), .A2(images_bus[425]), .A3(n8692), .ZN(n11829) );
  nd12d1 U8527 ( .A1(n6459), .A2(n3060), .ZN(n4733) );
  an02d1 U8532 ( .A1(N14274), .A2(n8691), .Z(n7939) );
  nr03d1 U8571 ( .A1(n11047), .A2(images_bus[433]), .A3(n3116), .ZN(n11836) );
  nr04d1 U8576 ( .A1(n6564), .A2(n7963), .A3(n3114), .A4(images_bus[435]), 
        .ZN(n11837) );
  nr03d1 U8601 ( .A1(n3011), .A2(images_bus[447]), .A3(n7973), .ZN(n5627) );
  an02d1 U8611 ( .A1(n2940), .A2(n11208), .Z(n4786) );
  nr03d1 U8612 ( .A1(n11853), .A2(n11852), .A3(n8031), .ZN(n11208) );
  an02d1 U8617 ( .A1(N14690), .A2(n3008), .Z(n9502) );
  nd04d1 U8635 ( .A1(n3005), .A2(n8047), .A3(n11860), .A4(n5979), .ZN(n11859)
         );
  nr03d1 U8658 ( .A1(n2966), .A2(images_bus[465]), .A3(n10369), .ZN(n7982) );
  nd12d1 U8669 ( .A1(n10258), .A2(n11877), .ZN(n10260) );
  nr03d1 U8673 ( .A1(n10362), .A2(images_bus[469]), .A3(n2973), .ZN(n11881) );
  nr03d1 U8681 ( .A1(n2980), .A2(images_bus[473]), .A3(n9538), .ZN(n11887) );
  nd04d1 U8683 ( .A1(n2979), .A2(n2977), .A3(n10357), .A4(n4890), .ZN(n11888)
         );
  nd04d1 U8695 ( .A1(n2828), .A2(n2842), .A3(n8796), .A4(n6074), .ZN(n11894)
         );
  an02d1 U8701 ( .A1(n4857), .A2(n4931), .Z(n5675) );
  an02d1 U8708 ( .A1(N15106), .A2(n11898), .Z(n10359) );
  nd04d1 U8717 ( .A1(n2913), .A2(n11126), .A3(n2852), .A4(n5221), .ZN(n11904)
         );
  nd04d1 U8731 ( .A1(n2877), .A2(n2876), .A3(n11187), .A4(n4393), .ZN(n11923)
         );
  nr04d1 U8735 ( .A1(images_bus[495]), .A2(n2909), .A3(n8810), .A4(n11186), 
        .ZN(n11925) );
  nr03d1 U8741 ( .A1(n11186), .A2(n2878), .A3(n2875), .ZN(n11919) );
  nr03d1 U8764 ( .A1(n2906), .A2(images_bus[499]), .A3(n11155), .ZN(n8013) );
  nd12d1 U8768 ( .A1(n4920), .A2(n11937), .ZN(n8008) );
  nr04d1 U8772 ( .A1(images_bus[503]), .A2(n10329), .A3(n9578), .A4(n2891), 
        .ZN(n11943) );
  an02d1 U8779 ( .A1(n2899), .A2(n11948), .Z(n11949) );
  an02d1 U8793 ( .A1(N15618), .A2(n11951), .Z(n11181) );
  an04d1 U8795 ( .A1(images_bus[509]), .A2(N15633), .A3(n11951), .A4(n12162), 
        .Z(n10341) );
  nd12d1 U8804 ( .A1(n9579), .A2(n8018), .ZN(n4916) );
  an03d1 U8810 ( .A1(n2894), .A2(n11953), .A3(N15554), .Z(n11175) );
  an02d1 U8813 ( .A1(images_bus[504]), .A2(n10329), .Z(n11953) );
  nr03d1 U8821 ( .A1(n6209), .A2(n9574), .A3(n5797), .ZN(n10329) );
  nr03d1 U8861 ( .A1(n6276), .A2(n11187), .A3(n5894), .ZN(n11931) );
  an02d1 U8887 ( .A1(N15298), .A2(n8798), .Z(n11190) );
  nd12d1 U8889 ( .A1(n10297), .A2(N15314), .ZN(n10307) );
  an03d1 U8897 ( .A1(images_bus[484]), .A2(images_bus[483]), .A3(n7341), .Z(
        n4926) );
  an02d1 U8905 ( .A1(n11965), .A2(n11193), .Z(n8802) );
  an02d1 U8906 ( .A1(n4869), .A2(n2859), .Z(n11193) );
  nr03d1 U8908 ( .A1(n10296), .A2(images_bus[487]), .A3(n11191), .ZN(n11964)
         );
  nr03d1 U8910 ( .A1(n6356), .A2(n11130), .A3(n11960), .ZN(n8798) );
  an04d1 U8916 ( .A1(images_bus[487]), .A2(images_bus[486]), .A3(N15282), .A4(
        n2864), .Z(n11191) );
  an02d1 U8925 ( .A1(n2850), .A2(n5678), .Z(n5679) );
  an02d1 U8935 ( .A1(n7345), .A2(n6079), .Z(n4927) );
  an02d1 U8940 ( .A1(n8782), .A2(n7999), .Z(n11893) );
  nd12d1 U8952 ( .A1(n10282), .A2(N15202), .ZN(n10285) );
  an02d1 U8954 ( .A1(N15218), .A2(n10288), .Z(n4869) );
  nr03d1 U8958 ( .A1(n11903), .A2(n10280), .A3(n5715), .ZN(n8831) );
  an02d1 U8961 ( .A1(n8783), .A2(n6425), .Z(n11898) );
  nr03d1 U8974 ( .A1(n6655), .A2(n11966), .A3(n4890), .ZN(n8783) );
  an02d1 U8979 ( .A1(n7989), .A2(n4299), .Z(n4936) );
  nd12d1 U9006 ( .A1(n7332), .A2(N15010), .ZN(n7333) );
  nd12d1 U9009 ( .A1(n10362), .A2(n2973), .ZN(n4839) );
  nr03d1 U9019 ( .A1(n7985), .A2(n11878), .A3(n4820), .ZN(n4938) );
  an02d1 U9051 ( .A1(n11861), .A2(n4940), .Z(n11868) );
  an02d1 U9052 ( .A1(n7317), .A2(n7360), .Z(n4940) );
  an03d1 U9053 ( .A1(images_bus[456]), .A2(images_bus[455]), .A3(n9510), .Z(
        n7360) );
  nd12d1 U9069 ( .A1(n10240), .A2(N14866), .ZN(n7359) );
  nr03d1 U9095 ( .A1(n5979), .A2(n10230), .A3(n7117), .ZN(n7311) );
  an02d1 U9109 ( .A1(N14754), .A2(n2951), .Z(n8047) );
  an03d1 U9138 ( .A1(n3013), .A2(n11854), .A3(images_bus[447]), .Z(n8738) );
  nr04d1 U9174 ( .A1(images_bus[443]), .A2(n3104), .A3(n6557), .A4(n11071), 
        .ZN(n11977) );
  an02d1 U9191 ( .A1(n6561), .A2(n3112), .Z(n10203) );
  an02d1 U9224 ( .A1(N14434), .A2(n3115), .Z(n9601) );
  an03d1 U9247 ( .A1(n5621), .A2(n8691), .A3(images_bus[427]), .Z(n6456) );
  an02d1 U9252 ( .A1(images_bus[421]), .A2(n6442), .Z(n9459) );
  an02d1 U9258 ( .A1(n10172), .A2(n6599), .Z(n6442) );
  an02d1 U9276 ( .A1(N14146), .A2(n3044), .Z(n7922) );
  an03d1 U9291 ( .A1(images_bus[414]), .A2(n6430), .A3(images_bus[415]), .Z(
        n11981) );
  nr03d1 U9315 ( .A1(n5709), .A2(n5552), .A3(n4900), .ZN(n8670) );
  nr03d1 U9324 ( .A1(n8057), .A2(n3222), .A3(n3213), .ZN(n5554) );
  nd12d1 U9359 ( .A1(n9436), .A2(N13922), .ZN(n8836) );
  an02d1 U9375 ( .A1(n8635), .A2(n11986), .Z(n5537) );
  an03d1 U9402 ( .A1(images_bus[395]), .A2(n11989), .A3(images_bus[396]), .Z(
        n9429) );
  nr03d1 U9405 ( .A1(n6558), .A2(n5145), .A3(n6591), .ZN(n5712) );
  an02d1 U9419 ( .A1(N13762), .A2(n6373), .Z(n9425) );
  an02d1 U9432 ( .A1(images_bus[394]), .A2(n11992), .Z(n11989) );
  an02d1 U9434 ( .A1(images_bus[393]), .A2(n6373), .Z(n11992) );
  an02d1 U9435 ( .A1(images_bus[392]), .A2(n11991), .Z(n6373) );
  an02d1 U9436 ( .A1(images_bus[391]), .A2(n8624), .Z(n11991) );
  an03d1 U9447 ( .A1(images_bus[389]), .A2(n4645), .A3(images_bus[390]), .Z(
        n4967) );
  an02d1 U9449 ( .A1(n11782), .A2(n4968), .Z(n11993) );
  nr03d1 U9452 ( .A1(n4969), .A2(n4970), .A3(n11774), .ZN(n11782) );
  nd12d1 U9480 ( .A1(n9422), .A2(N13714), .ZN(n6378) );
  nd12d1 U9488 ( .A1(n7215), .A2(images_bus[385]), .ZN(n6363) );
  nr03d1 U9490 ( .A1(n6162), .A2(n7209), .A3(n6089), .ZN(n11779) );
  an02d1 U9499 ( .A1(images_bus[380]), .A2(n6340), .Z(n10958) );
  an02d1 U9503 ( .A1(images_bus[379]), .A2(n8838), .Z(n6340) );
  an02d1 U9504 ( .A1(n10109), .A2(n6664), .Z(n8838) );
  an02d1 U9506 ( .A1(images_bus[377]), .A2(n5718), .Z(n10109) );
  an02d1 U9511 ( .A1(N13426), .A2(n7190), .Z(n7189) );
  nd12d1 U9521 ( .A1(n5504), .A2(N13458), .ZN(n5501) );
  an02d1 U9525 ( .A1(images_bus[372]), .A2(n7190), .Z(n8601) );
  an02d1 U9526 ( .A1(images_bus[371]), .A2(n10099), .Z(n7190) );
  an02d1 U9534 ( .A1(n5488), .A2(n6737), .Z(n10099) );
  an02d1 U9538 ( .A1(N13378), .A2(n8069), .Z(n10935) );
  an02d1 U9541 ( .A1(images_bus[369]), .A2(n8069), .Z(n5488) );
  nr03d1 U9549 ( .A1(n6318), .A2(n4611), .A3(n6597), .ZN(n5717) );
  nd12d1 U9564 ( .A1(n11743), .A2(n4977), .ZN(n11746) );
  nr03d1 U9572 ( .A1(n4979), .A2(n4591), .A3(n11733), .ZN(n11736) );
  nd12d1 U9575 ( .A1(n7381), .A2(n11752), .ZN(n4602) );
  an02d1 U9585 ( .A1(n11748), .A2(n7169), .Z(n11999) );
  nd12d1 U9587 ( .A1(n5485), .A2(N13282), .ZN(n7381) );
  an02d1 U9592 ( .A1(n12000), .A2(n5626), .Z(n7384) );
  an02d1 U9595 ( .A1(images_bus[360]), .A2(n10918), .Z(n12000) );
  an02d1 U9600 ( .A1(n11741), .A2(n6601), .Z(n7160) );
  an04d1 U9611 ( .A1(n3275), .A2(n3273), .A3(n3330), .A4(n12001), .Z(n4582) );
  nd12d1 U9624 ( .A1(n7147), .A2(N13106), .ZN(n5474) );
  nr03d1 U9626 ( .A1(n4982), .A2(n4981), .A3(n11719), .ZN(n11731) );
  nd12d1 U9627 ( .A1(n11715), .A2(n4983), .ZN(n11719) );
  an02d1 U9628 ( .A1(n6243), .A2(n5723), .Z(n4983) );
  an02d1 U9651 ( .A1(images_bus[349]), .A2(n5463), .Z(n6271) );
  nr03d1 U9655 ( .A1(n11729), .A2(n5463), .A3(n3391), .ZN(n4570) );
  nd12d1 U9659 ( .A1(n8572), .A2(N13042), .ZN(n8579) );
  an02d1 U9672 ( .A1(images_bus[345]), .A2(n12005), .Z(n12004) );
  an02d1 U9673 ( .A1(images_bus[344]), .A2(n11723), .Z(n12005) );
  an02d1 U9674 ( .A1(images_bus[343]), .A2(n11726), .Z(n11723) );
  nd12d1 U9687 ( .A1(n11716), .A2(N12898), .ZN(n6252) );
  nr04d1 U9697 ( .A1(n9342), .A2(n6241), .A3(n7132), .A4(n12008), .ZN(n4986)
         );
  an03d1 U9704 ( .A1(images_bus[336]), .A2(n12010), .A3(images_bus[337]), .Z(
        n12007) );
  an03d1 U9705 ( .A1(images_bus[336]), .A2(n12010), .A3(N12866), .Z(n7128) );
  an02d1 U9706 ( .A1(n11703), .A2(n4988), .Z(n11711) );
  an02d1 U9707 ( .A1(n5725), .A2(n5634), .Z(n4988) );
  an02d1 U9723 ( .A1(N12850), .A2(n12010), .Z(n10882) );
  an02d1 U9726 ( .A1(images_bus[333]), .A2(n9610), .Z(n12012) );
  an02d1 U9727 ( .A1(images_bus[332]), .A2(n12009), .Z(n9610) );
  an02d1 U9728 ( .A1(images_bus[331]), .A2(n11709), .Z(n12009) );
  an02d1 U9729 ( .A1(images_bus[330]), .A2(n8852), .Z(n11709) );
  an02d1 U9730 ( .A1(images_bus[329]), .A2(n11710), .Z(n8852) );
  an02d1 U9731 ( .A1(images_bus[328]), .A2(n12015), .Z(n11710) );
  nr03d1 U9737 ( .A1(n4990), .A2(n4989), .A3(n11705), .ZN(n11703) );
  nd12d1 U9745 ( .A1(n10861), .A2(N12674), .ZN(n10863) );
  an02d1 U9754 ( .A1(images_bus[327]), .A2(n12017), .Z(n12015) );
  an02d1 U9763 ( .A1(images_bus[323]), .A2(n11697), .Z(n11696) );
  an02d1 U9764 ( .A1(images_bus[322]), .A2(n10054), .Z(n11697) );
  an02d1 U9767 ( .A1(images_bus[323]), .A2(n6603), .Z(n4537) );
  an02d1 U9776 ( .A1(images_bus[321]), .A2(n5422), .Z(n10054) );
  an02d1 U9777 ( .A1(images_bus[320]), .A2(n12018), .Z(n5422) );
  nr03d1 U9780 ( .A1(n4526), .A2(n6098), .A3(n7232), .ZN(n4991) );
  nr03d1 U9783 ( .A1(n4993), .A2(n4992), .A3(n11685), .ZN(n11687) );
  an02d1 U9785 ( .A1(n5731), .A2(n11677), .Z(n4994) );
  nr03d1 U9808 ( .A1(n10847), .A2(images_bus[315]), .A3(n9315), .ZN(n7807) );
  an02d1 U9816 ( .A1(images_bus[313]), .A2(n6193), .Z(n11680) );
  an02d1 U9817 ( .A1(n5833), .A2(n10837), .Z(n6193) );
  an02d1 U9820 ( .A1(n5052), .A2(n11681), .Z(n11679) );
  nd04d1 U9838 ( .A1(images_bus[305]), .A2(N12370), .A3(images_bus[304]), .A4(
        n3439), .ZN(n7085) );
  an03d1 U9841 ( .A1(N12354), .A2(n3439), .A3(images_bus[304]), .Z(n11673) );
  nr03d1 U9846 ( .A1(n5398), .A2(n6608), .A3(n8518), .ZN(n4996) );
  an03d1 U9847 ( .A1(n6018), .A2(n4677), .A3(n12021), .Z(n4492) );
  an03d1 U9858 ( .A1(N12306), .A2(n3461), .A3(images_bus[301]), .Z(n11668) );
  an03d1 U9872 ( .A1(n3467), .A2(n5642), .A3(N12258), .Z(n10825) );
  nr03d1 U9875 ( .A1(n10823), .A2(n8518), .A3(n5396), .ZN(n12022) );
  an02d1 U9881 ( .A1(n4677), .A2(n5384), .Z(n7064) );
  nd12d1 U9890 ( .A1(n6172), .A2(N12146), .ZN(n6169) );
  an03d1 U9912 ( .A1(images_bus[287]), .A2(n7046), .A3(images_bus[288]), .Z(
        n4484) );
  an03d1 U9916 ( .A1(N12082), .A2(n7046), .A3(images_bus[287]), .Z(n9276) );
  an02d1 U9917 ( .A1(images_bus[286]), .A2(n5377), .Z(n7046) );
  nr03d1 U9918 ( .A1(n12026), .A2(n12149), .A3(n3478), .ZN(n5377) );
  an03d1 U9920 ( .A1(n5000), .A2(images_bus[288]), .A3(n3508), .Z(n11656) );
  nr03d1 U9935 ( .A1(n7016), .A2(n9620), .A3(n5741), .ZN(n5001) );
  an02d1 U9942 ( .A1(n12027), .A2(n12028), .Z(n4461) );
  nd04d1 U9945 ( .A1(images_bus[281]), .A2(N11986), .A3(images_bus[280]), .A4(
        n12032), .ZN(n6151) );
  an02d1 U9951 ( .A1(n5413), .A2(n12032), .Z(n10795) );
  an02d1 U9956 ( .A1(n6148), .A2(n3543), .Z(n4468) );
  an02d1 U9959 ( .A1(N11954), .A2(n12032), .Z(n10788) );
  nd12d1 U9984 ( .A1(n11642), .A2(n5002), .ZN(n11645) );
  an02d1 U9991 ( .A1(N11858), .A2(n5362), .Z(n9998) );
  an02d1 U9996 ( .A1(n6614), .A2(n3563), .Z(n5362) );
  an02d1 U9997 ( .A1(images_bus[273]), .A2(n5002), .Z(n6614) );
  an03d1 U10002 ( .A1(n5002), .A2(n3563), .A3(N11842), .Z(n7040) );
  nd12d1 U10009 ( .A1(n8482), .A2(n9246), .ZN(n8076) );
  an03d1 U10016 ( .A1(N11794), .A2(n12040), .A3(images_bus[269]), .Z(n10400)
         );
  nd04d1 U10028 ( .A1(n5647), .A2(n9248), .A3(images_bus[264]), .A4(n8477), 
        .ZN(n5005) );
  an02d1 U10041 ( .A1(images_bus[268]), .A2(n12041), .Z(n12040) );
  an03d1 U10042 ( .A1(images_bus[266]), .A2(n9977), .A3(images_bus[267]), .Z(
        n12041) );
  an03d1 U10064 ( .A1(n12047), .A2(images_bus[262]), .A3(N11682), .Z(n8471) );
  an02d1 U10067 ( .A1(n10402), .A2(n8855), .Z(n12047) );
  an02d1 U10068 ( .A1(images_bus[259]), .A2(n9621), .Z(n8855) );
  nr03d1 U10072 ( .A1(n5746), .A2(n11253), .A3(n6923), .ZN(n10402) );
  nr03d1 U10082 ( .A1(n11610), .A2(n5750), .A3(n12048), .ZN(n11625) );
  an03d1 U10106 ( .A1(n3787), .A2(images_bus[249]), .A3(N11481), .Z(n5337) );
  nd12d1 U10123 ( .A1(n9222), .A2(n9223), .ZN(n7002) );
  an03d1 U10124 ( .A1(N11421), .A2(n3798), .A3(images_bus[245]), .Z(n9223) );
  an02d1 U10146 ( .A1(n5752), .A2(n5303), .Z(n6087) );
  an02d1 U10181 ( .A1(n6976), .A2(n6621), .Z(n9199) );
  nr03d1 U10185 ( .A1(n7242), .A2(n11586), .A3(n5747), .ZN(n8433) );
  nd12d1 U10197 ( .A1(n11576), .A2(n5759), .ZN(n11579) );
  an02d1 U10202 ( .A1(n5758), .A2(n5433), .Z(n6623) );
  nr03d1 U10204 ( .A1(n7019), .A2(n5839), .A3(n7704), .ZN(n5758) );
  nd12d1 U10208 ( .A1(n5270), .A2(n3736), .ZN(n9935) );
  nd12d1 U10225 ( .A1(n5248), .A2(n5240), .ZN(n7418) );
  an02d1 U10228 ( .A1(N10941), .A2(n3870), .Z(n5240) );
  an03d1 U10238 ( .A1(images_bus[208]), .A2(images_bus[207]), .A3(n8864), .Z(
        n6624) );
  nr03d1 U10239 ( .A1(n6571), .A2(n5186), .A3(n5218), .ZN(n8864) );
  nd12d1 U10245 ( .A1(n10688), .A2(N10821), .ZN(n7690) );
  an02d1 U10252 ( .A1(n7696), .A2(n7697), .Z(n7691) );
  an03d1 U10253 ( .A1(n5232), .A2(n3874), .A3(n3875), .Z(n7696) );
  an02d1 U10254 ( .A1(N10896), .A2(n3873), .Z(n5232) );
  nr03d1 U10276 ( .A1(n5225), .A2(n9911), .A3(n5227), .ZN(n7697) );
  nr03d1 U10283 ( .A1(n5209), .A2(n12128), .A3(n5186), .ZN(n9167) );
  nd12d1 U10286 ( .A1(n8400), .A2(n7685), .ZN(n5210) );
  nr03d1 U10305 ( .A1(n5276), .A2(n9903), .A3(n6628), .ZN(n5201) );
  nd12d1 U10307 ( .A1(n11565), .A2(n5765), .ZN(n11568) );
  an03d1 U10319 ( .A1(images_bus[195]), .A2(n3835), .A3(N10671), .Z(n10676) );
  an02d1 U10330 ( .A1(n4957), .A2(n5767), .Z(n7423) );
  an02d1 U10333 ( .A1(N10611), .A2(n3828), .Z(n5770) );
  nr03d1 U10368 ( .A1(n6921), .A2(n6631), .A3(n5774), .ZN(n5181) );
  nr03d1 U10377 ( .A1(n7427), .A2(n8373), .A3(n4316), .ZN(n9139) );
  an02d1 U10395 ( .A1(n6906), .A2(n3935), .Z(n5163) );
  an03d1 U10398 ( .A1(images_bus[175]), .A2(n9876), .A3(N10371), .Z(n6906) );
  an02d1 U10399 ( .A1(n4470), .A2(n6902), .Z(n9876) );
  nr04d1 U10404 ( .A1(n11524), .A2(n5139), .A3(n8093), .A4(n7433), .ZN(n11536)
         );
  nr03d1 U10413 ( .A1(n10640), .A2(n4464), .A3(n4422), .ZN(n8361) );
  nd04d1 U10417 ( .A1(N10281), .A2(n3963), .A3(images_bus[168]), .A4(
        images_bus[169]), .ZN(n6896) );
  an03d1 U10422 ( .A1(n3930), .A2(images_bus[171]), .A3(N10311), .Z(n11534) );
  an02d1 U10444 ( .A1(N10146), .A2(n9857), .Z(n5120) );
  an03d1 U10445 ( .A1(images_bus[159]), .A2(n7648), .A3(images_bus[160]), .Z(
        n9857) );
  an02d1 U10453 ( .A1(n11519), .A2(images_bus[159]), .Z(n11517) );
  nr04d1 U10454 ( .A1(n11508), .A2(n5112), .A3(n7640), .A4(n7645), .ZN(n11519)
         );
  nr03d1 U10460 ( .A1(n7023), .A2(n5099), .A3(n5440), .ZN(n8340) );
  an02d1 U10468 ( .A1(N10011), .A2(n4037), .Z(n10617) );
  an02d1 U10471 ( .A1(n8095), .A2(n11271), .Z(n7633) );
  an03d1 U10472 ( .A1(images_bus[150]), .A2(n4048), .A3(N9996), .Z(n11271) );
  an02d1 U10474 ( .A1(N9966), .A2(n4047), .Z(n8095) );
  nr03d1 U10511 ( .A1(n5194), .A2(n11493), .A3(n6575), .ZN(n9104) );
  an03d1 U10515 ( .A1(n8870), .A2(n5687), .A3(n11487), .Z(n11491) );
  an02d1 U10527 ( .A1(images_bus[135]), .A2(n8317), .Z(n6851) );
  an03d1 U10529 ( .A1(images_bus[136]), .A2(images_bus[133]), .A3(n11480), .Z(
        n11487) );
  an02d1 U10531 ( .A1(N9756), .A2(n8317), .Z(n9098) );
  an02d1 U10541 ( .A1(n11482), .A2(images_bus[132]), .Z(n11480) );
  nr04d1 U10542 ( .A1(n3994), .A2(n5281), .A3(n6946), .A4(n5768), .ZN(n11482)
         );
  nr04d1 U10547 ( .A1(n11468), .A2(n9640), .A3(n7245), .A4(n6650), .ZN(n11478)
         );
  an02d1 U10575 ( .A1(N9582), .A2(n9081), .Z(n8876) );
  an02d1 U10579 ( .A1(n9081), .A2(images_bus[123]), .Z(n11470) );
  an02d1 U10603 ( .A1(n11431), .A2(n5890), .Z(n11435) );
  nr03d1 U10626 ( .A1(n5957), .A2(n4105), .A3(n7097), .ZN(n12065) );
  an03d1 U10638 ( .A1(images_bus[106]), .A2(n6790), .A3(images_bus[107]), .Z(
        n5911) );
  an03d1 U10644 ( .A1(images_bus[104]), .A2(n8282), .A3(images_bus[105]), .Z(
        n6790) );
  an02d1 U10653 ( .A1(N9274), .A2(n4113), .Z(n5895) );
  nd12d1 U10669 ( .A1(n7572), .A2(N9218), .ZN(n6781) );
  nr03d1 U10671 ( .A1(n4139), .A2(n7251), .A3(n11427), .ZN(n11431) );
  nd12d1 U10672 ( .A1(n11422), .A2(n6660), .ZN(n11427) );
  nd12d1 U10700 ( .A1(n5876), .A2(N9162), .ZN(n5027) );
  nr03d1 U10703 ( .A1(n7561), .A2(n7447), .A3(n4973), .ZN(n8268) );
  an03d1 U10709 ( .A1(images_bus[86]), .A2(n11286), .A3(images_bus[87]), .Z(
        n11423) );
  nr03d1 U10711 ( .A1(n6768), .A2(n11287), .A3(n5016), .ZN(n7557) );
  an03d1 U10713 ( .A1(images_bus[84]), .A2(n11416), .A3(images_bus[85]), .Z(
        n11286) );
  an02d1 U10721 ( .A1(n11417), .A2(images_bus[84]), .Z(n11419) );
  nr03d1 U10722 ( .A1(n6662), .A2(n5106), .A3(n11411), .ZN(n11417) );
  nd12d1 U10723 ( .A1(n5844), .A2(n11404), .ZN(n11411) );
  an02d1 U10727 ( .A1(n7548), .A2(n10542), .Z(n6762) );
  an03d1 U10728 ( .A1(n4179), .A2(n7450), .A3(N8994), .Z(n10542) );
  an03d1 U10747 ( .A1(n6663), .A2(images_bus[74]), .A3(n4145), .Z(n11404) );
  an02d1 U10761 ( .A1(N8882), .A2(n4182), .Z(n5828) );
  an02d1 U10767 ( .A1(N8840), .A2(n4184), .Z(n9008) );
  nr03d1 U10772 ( .A1(n6748), .A2(n4751), .A3(n11394), .ZN(n11395) );
  nd04d1 U10773 ( .A1(n5778), .A2(n4205), .A3(images_bus[67]), .A4(n12069), 
        .ZN(n11394) );
  an03d1 U10814 ( .A1(images_bus[44]), .A2(images_bus[43]), .A3(n11355), .Z(
        n11356) );
  an02d1 U10817 ( .A1(n8118), .A2(images_bus[48]), .Z(n7456) );
  an02d1 U10832 ( .A1(images_bus[56]), .A2(n11375), .Z(n12071) );
  nr03d1 U10833 ( .A1(n6270), .A2(n11373), .A3(n5862), .ZN(n11375) );
  an03d1 U10838 ( .A1(n8197), .A2(n6719), .A3(images_bus[48]), .Z(n6720) );
  nd12d1 U10851 ( .A1(n8195), .A2(n11357), .ZN(n5800) );
  nd12d1 U10853 ( .A1(n10491), .A2(N8510), .ZN(n8195) );
  an02d1 U10866 ( .A1(images_bus[41]), .A2(n8188), .Z(n10426) );
  an02d1 U10867 ( .A1(n4275), .A2(n6702), .Z(n8188) );
  an02d1 U10878 ( .A1(n11344), .A2(n6697), .Z(n11346) );
  nd04d1 U10894 ( .A1(N8393), .A2(N8380), .A3(n9697), .A4(images_bus[35]), 
        .ZN(n8937) );
  an02d1 U10895 ( .A1(n11342), .A2(n6967), .Z(n9697) );
  nd12d1 U10897 ( .A1(n10478), .A2(n11342), .ZN(n6686) );
  an02d1 U10919 ( .A1(N8318), .A2(n10468), .Z(n8174) );
  an02d1 U10920 ( .A1(N8306), .A2(n11336), .Z(n10468) );
  an02d1 U10923 ( .A1(images_bus[27]), .A2(n7487), .Z(n8127) );
  nd12d1 U10927 ( .A1(n8165), .A2(n8161), .ZN(n9684) );
  an02d1 U10931 ( .A1(N8258), .A2(n11333), .Z(n8161) );
  nd12d1 U10935 ( .A1(n11330), .A2(N8246), .ZN(n7485) );
  nr03d1 U10949 ( .A1(n4608), .A2(n10445), .A3(n6355), .ZN(n8147) );
  an03d1 U10975 ( .A1(n11304), .A2(images_bus[4]), .A3(N8034), .Z(n8894) );
  nr03d1 U10976 ( .A1(n6975), .A2(n5785), .A3(n5315), .ZN(n11304) );
  reordering_DW01_inc_0_DW01_inc_2 add_174 ( .A({count_image[8:6], 
        \lt_82/A[5] , \lt_82/A[4] , count_image[3:0]}), .SUM({N6845, N6844, 
        N6843, N6842, N6841, N6840, N6839, N6838, N6837}) );
  reordering_DW01_add_9 add_0_root_add_86_root_add_255_countones_143 ( .A({
        1'b0, 1'b0, N28504, N28503, N28502, N28501, N28500, N28499, N28498}), 
        .B({1'b0, N28613, N28612, N28611, N28610, N28609, N28608, N28607, 
        N28606}), .CI(1'b0), .SUM({N5028, N5027, N5026, N5025, N5024, N5023, 
        N5022, N5021, N5020}) );
  reordering_DW01_inc_1_DW01_inc_6 r7602 ( .A({n510, N3181, n508, n506, n504, 
        n955, N3974, n500, n513}), .SUM({N4013, N4012, N4011, N4010, N5074, 
        N5073, N5072, N5071, N5070}) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28355), .B(
        N28571), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_1_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28607) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28356), .B(
        N28572), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_1_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28608) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28357), .B(
        N28573), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_1_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28609) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_4  ( .A(N28358), .B(
        N28574), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(\add_1_root_add_86_root_add_255_countones_143/carry[5] ), .S(
        N28610) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_5  ( .A(N28359), .B(
        N28575), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[5] ), 
        .CO(\add_1_root_add_86_root_add_255_countones_143/carry[6] ), .S(
        N28611) );
  ad01d0 \add_1_root_add_86_root_add_255_countones_143/U1_6  ( .A(N28360), .B(
        N28576), .CI(\add_1_root_add_86_root_add_255_countones_143/carry[6] ), 
        .CO(N28613), .S(N28612) );
  ad01d0 \add_2_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27491), .B(
        N28076), .CI(\add_2_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_2_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28571) );
  ad01d0 \add_2_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27492), .B(
        N28077), .CI(\add_2_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_2_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28572) );
  ad01d0 \add_2_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27493), .B(
        N28078), .CI(\add_2_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_2_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28573) );
  ad01d0 \add_2_root_add_86_root_add_255_countones_143/U1_4  ( .A(N27494), .B(
        N28079), .CI(\add_2_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(\add_2_root_add_86_root_add_255_countones_143/carry[5] ), .S(
        N28574) );
  ad01d0 \add_2_root_add_86_root_add_255_countones_143/U1_5  ( .A(N27495), .B(
        N28080), .CI(\add_2_root_add_86_root_add_255_countones_143/carry[5] ), 
        .CO(N28576), .S(N28575) );
  ad01d0 \add_3_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27500), .B(
        N28067), .CI(\add_3_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_3_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28499) );
  ad01d0 \add_3_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27501), .B(
        N28068), .CI(\add_3_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_3_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28500) );
  ad01d0 \add_3_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27502), .B(
        N28069), .CI(\add_3_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_3_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28501) );
  ad01d0 \add_3_root_add_86_root_add_255_countones_143/U1_4  ( .A(N27503), .B(
        N28070), .CI(\add_3_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(\add_3_root_add_86_root_add_255_countones_143/carry[5] ), .S(
        N28502) );
  ad01d0 \add_3_root_add_86_root_add_255_countones_143/U1_5  ( .A(N27504), .B(
        N28071), .CI(\add_3_root_add_86_root_add_255_countones_143/carry[5] ), 
        .CO(N28504), .S(N28503) );
  ad01d0 \add_4_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28364), .B(
        N27509), .CI(\add_4_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_4_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28355) );
  ad01d0 \add_4_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28365), .B(
        N27510), .CI(\add_4_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_4_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28356) );
  ad01d0 \add_4_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28366), .B(
        N27511), .CI(\add_4_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_4_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28357) );
  ad01d0 \add_4_root_add_86_root_add_255_countones_143/U1_4  ( .A(N28367), .B(
        N27512), .CI(\add_4_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(\add_4_root_add_86_root_add_255_countones_143/carry[5] ), .S(
        N28358) );
  ad01d0 \add_11_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27590), 
        .B(N27581), .CI(
        \add_11_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_11_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28364)
         );
  ad01d0 \add_11_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27591), 
        .B(N27582), .CI(
        \add_11_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_11_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28365)
         );
  ad01d0 \add_11_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27592), 
        .B(N27583), .CI(
        \add_11_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N28367), 
        .S(N28366) );
  ad01d0 \add_8_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28373), .B(
        N28508), .CI(\add_8_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_8_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28076) );
  ad01d0 \add_8_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28374), .B(
        N28509), .CI(\add_8_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_8_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28077) );
  ad01d0 \add_8_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28375), .B(
        N28510), .CI(\add_8_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_8_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28078) );
  ad01d0 \add_8_root_add_86_root_add_255_countones_143/U1_4  ( .A(N28376), .B(
        N28511), .CI(\add_8_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(N28080), .S(N28079) );
  ad01d0 \add_18_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27644), 
        .B(N28121), .CI(
        \add_18_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_18_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28508)
         );
  ad01d0 \add_18_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27645), 
        .B(N28122), .CI(
        \add_18_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_18_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28509)
         );
  ad01d0 \add_18_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27646), 
        .B(N28123), .CI(
        \add_18_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N28511), 
        .S(N28510) );
  ad01d0 \add_27_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28193), 
        .B(N27689), .CI(
        \add_27_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_27_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28121)
         );
  ad01d0 \add_27_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28194), 
        .B(N27690), .CI(
        \add_27_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28123), 
        .S(N28122) );
  ad01d0 \add_58_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27968), 
        .B(N27455), .CI(
        \add_58_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28194), 
        .S(N28193) );
  ad01d0 \add_19_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27635), 
        .B(N27563), .CI(
        \add_19_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_19_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28373)
         );
  ad01d0 \add_19_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27636), 
        .B(N27564), .CI(
        \add_19_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_19_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28374)
         );
  ad01d0 \add_19_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27637), 
        .B(N27565), .CI(
        \add_19_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N28376), 
        .S(N28375) );
  ad01d0 \add_5_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28085), .B(
        N27554), .CI(\add_5_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_5_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N28067) );
  ad01d0 \add_5_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28086), .B(
        N27555), .CI(\add_5_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_5_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N28068) );
  ad01d0 \add_5_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28087), .B(
        N27556), .CI(\add_5_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_5_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N28069) );
  ad01d0 \add_5_root_add_86_root_add_255_countones_143/U1_4  ( .A(N28088), .B(
        N27557), .CI(\add_5_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(N28071), .S(N28070) );
  ad01d0 \add_12_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28382), 
        .B(N27599), .CI(
        \add_12_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_12_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28085)
         );
  ad01d0 \add_12_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28383), 
        .B(N27600), .CI(
        \add_12_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_12_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28086)
         );
  ad01d0 \add_12_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28384), 
        .B(N27601), .CI(
        \add_12_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N28088), 
        .S(N28087) );
  ad01d0 \add_26_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28526), 
        .B(N28184), .CI(
        \add_26_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_26_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28382)
         );
  ad01d0 \add_26_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28527), 
        .B(N28185), .CI(
        \add_26_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28384), 
        .S(N28383) );
  ad01d0 \add_54_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28346), 
        .B(N27131), .CI(
        \add_54_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28185), 
        .S(N28184) );
  ad01d0 \add_162_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4926), 
        .B(N4785), .CI(N4782), .CO(N28346), .S(N28345) );
  ad01d0 \add_49_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28265), 
        .B(N28454), .CI(
        \add_49_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28527), 
        .S(N28526) );
  ad01d0 \add_91_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5002), .B(
        N4828), .CI(N4777), .CO(N28454), .S(N28453) );
  ad01d0 \add_92_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4801), .B(
        N4822), .CI(N4948), .CO(N28265), .S(N28264) );
  ad01d0 \add_128_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4973), 
        .B(N4901), .CI(N4799), .CO(N27968), .S(N27967) );
  ad01d0 \add_47_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27977), 
        .B(N27914), .CI(
        \add_47_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27690), 
        .S(N27689) );
  ad01d0 \add_103_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4891), 
        .B(N4882), .CI(N5014), .CO(N27914), .S(N27913) );
  ad01d0 \add_132_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4967), 
        .B(N4790), .CI(N4787), .CO(N27977), .S(N27976) );
  ad01d0 \add_38_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27806), 
        .B(N28589), .CI(
        \add_38_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_38_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27644)
         );
  ad01d0 \add_38_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27807), 
        .B(N28590), .CI(
        \add_38_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27646), 
        .S(N27645) );
  ad01d0 \add_65_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27221), 
        .B(N27410), .CI(
        \add_65_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28590), 
        .S(N28589) );
  ad01d0 \add_73_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28058), 
        .B(N28013), .CI(
        \add_73_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27807), 
        .S(N27806) );
  ad01d0 \add_148_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4995), 
        .B(N4848), .CI(N4941), .CO(N28013), .S(N28012) );
  ad01d0 \add_166_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4764), 
        .B(N4767), .CI(N4887), .CO(N28058), .S(N28057) );
  ad01d0 \add_37_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27815), 
        .B(N28535), .CI(
        \add_37_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_37_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27635)
         );
  ad01d0 \add_37_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27816), 
        .B(N28536), .CI(
        \add_37_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27637), 
        .S(N27636) );
  ad01d0 \add_66_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27185), 
        .B(N27365), .CI(
        \add_66_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28536), 
        .S(N28535) );
  ad01d0 \add_76_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27356), 
        .B(N27212), .CI(
        \add_76_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27816), 
        .S(N27815) );
  ad01d0 \add_28_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27725), 
        .B(N28166), .CI(
        \add_28_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_28_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27599)
         );
  ad01d0 \add_28_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27726), 
        .B(N28167), .CI(
        \add_28_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27601), 
        .S(N27600) );
  ad01d0 \add_46_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27941), 
        .B(N27113), .CI(
        \add_46_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28167), 
        .S(N28166) );
  ad01d0 \add_117_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4847), 
        .B(N4997), .CI(N4994), .CO(N27941), .S(N27940) );
  ad01d0 \add_55_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27230), 
        .B(N28049), .CI(
        \add_55_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27726), 
        .S(N27725) );
  ad01d0 \add_163_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4962), 
        .B(N4779), .CI(N4776), .CO(N28049), .S(N28048) );
  ad01d0 \add_25_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27707), 
        .B(N27770), .CI(
        \add_25_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_25_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27590)
         );
  ad01d0 \add_25_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27708), 
        .B(N27771), .CI(
        \add_25_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27592), 
        .S(N27591) );
  ad01d0 \add_63_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27419), 
        .B(N27374), .CI(
        \add_63_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27771), 
        .S(N27770) );
  ad01d0 \add_52_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28040), 
        .B(N27248), .CI(
        \add_52_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27708), 
        .S(N27707) );
  ad01d0 \add_159_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4797), 
        .B(N4971), .CI(N4794), .CO(N28040), .S(N28039) );
  ad01d0 \add_24_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28175), 
        .B(N27734), .CI(
        \add_24_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_24_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27581)
         );
  ad01d0 \add_24_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28176), 
        .B(N27735), .CI(
        \add_24_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27583), 
        .S(N27582) );
  ad01d0 \add_56_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27932), 
        .B(N28301), .CI(
        \add_56_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27735), 
        .S(N27734) );
  ad01d0 \add_124_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4817), 
        .B(N4937), .CI(N4913), .CO(N28301), .S(N28300) );
  ad01d0 \add_113_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4877), 
        .B(N4940), .CI(N5009), .CO(N27932), .S(N27931) );
  ad01d0 \add_51_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28472), 
        .B(N27464), .CI(
        \add_51_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28176), 
        .S(N28175) );
  ad01d0 \add_123_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4982), 
        .B(N4823), .CI(N4820), .CO(N28472), .S(N28471) );
  ad01d0 \add_21_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27752), 
        .B(N28427), .CI(
        \add_21_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_21_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27563)
         );
  ad01d0 \add_21_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27753), 
        .B(N28428), .CI(
        \add_21_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27565), 
        .S(N27564) );
  ad01d0 \add_67_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27986), 
        .B(N28490), .CI(
        \add_67_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28428), 
        .S(N28427) );
  ad01d0 \add_154_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4899), 
        .B(N4911), .CI(N4893), .CO(N28490), .S(N28489) );
  ad01d0 \add_135_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4880), 
        .B(N4895), .CI(N4961), .CO(N27986), .S(N27985) );
  ad01d0 \add_60_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27428), 
        .B(N28328), .CI(
        \add_60_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27753), 
        .S(N27752) );
  ad01d0 \add_147_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4851), 
        .B(N4854), .CI(N4998), .CO(N28328), .S(N28327) );
  ad01d0 \add_17_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28139), 
        .B(N27626), .CI(
        \add_17_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_17_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27554)
         );
  ad01d0 \add_17_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28140), 
        .B(N27627), .CI(
        \add_17_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_17_root_add_86_root_add_255_countones_143/carry[3] ), .S(N27555)
         );
  ad01d0 \add_17_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28141), 
        .B(N27628), .CI(
        \add_17_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N27557), 
        .S(N27556) );
  ad01d0 \add_32_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27797), 
        .B(N27833), .CI(
        \add_32_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_32_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27626)
         );
  ad01d0 \add_32_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27798), 
        .B(N27834), .CI(
        \add_32_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27628), 
        .S(N27627) );
  ad01d0 \add_79_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27302), 
        .B(N28283), .CI(
        \add_79_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27834), 
        .S(N27833) );
  ad01d0 \add_109_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4765), 
        .B(N4906), .CI(N4921), .CO(N28283), .S(N28282) );
  ad01d0 \add_72_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28598), 
        .B(N28553), .CI(
        \add_72_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27798), 
        .S(N27797) );
  ad01d0 \add_107_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4888), 
        .B(N4924), .CI(N4957), .CO(N28553), .S(N28552) );
  ad01d0 \add_106_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4987), 
        .B(N4885), .CI(N4771), .CO(N28598), .S(N28597) );
  ad01d0 \add_36_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28229), 
        .B(N27842), .CI(
        \add_36_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_36_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28139)
         );
  ad01d0 \add_36_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28230), 
        .B(N27843), .CI(
        \add_36_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28141), 
        .S(N28140) );
  ad01d0 \add_80_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28031), 
        .B(N28562), .CI(
        \add_80_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27843), 
        .S(N27842) );
  ad01d0 \add_138_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4907), 
        .B(N4922), .CI(N4766), .CO(N28562), .S(N28561) );
  ad01d0 \add_156_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4812), 
        .B(N4980), .CI(N4809), .CO(N28031), .S(N28030) );
  ad01d0 \add_75_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27347), 
        .B(N27473), .CI(
        \add_75_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28230), 
        .S(N28229) );
  ad01d0 \add_9_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28103), .B(
        N27518), .CI(\add_9_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_9_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N27509) );
  ad01d0 \add_9_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28104), .B(
        N27519), .CI(\add_9_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_9_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N27510) );
  ad01d0 \add_9_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28105), .B(
        N27520), .CI(\add_9_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_9_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N27511) );
  ad01d0 \add_9_root_add_86_root_add_255_countones_143/U1_4  ( .A(N28106), .B(
        N27521), .CI(\add_9_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(N27513), .S(N27512) );
  ad01d0 \add_10_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27617), 
        .B(N28391), .CI(
        \add_10_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_10_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27518)
         );
  ad01d0 \add_10_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27618), 
        .B(N28392), .CI(
        \add_10_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_10_root_add_86_root_add_255_countones_143/carry[3] ), .S(N27519)
         );
  ad01d0 \add_10_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27619), 
        .B(N28393), .CI(
        \add_10_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N27521), 
        .S(N27520) );
  ad01d0 \add_35_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28220), 
        .B(N28211), .CI(
        \add_35_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_35_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28391)
         );
  ad01d0 \add_35_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28221), 
        .B(N28212), .CI(
        \add_35_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28393), 
        .S(N28392) );
  ad01d0 \add_68_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27482), 
        .B(N27167), .CI(
        \add_68_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28212), 
        .S(N28211) );
  ad01d0 \add_71_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28310), 
        .B(N28319), .CI(
        \add_71_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28221), 
        .S(N28220) );
  ad01d0 \add_140_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4884), 
        .B(N4946), .CI(N5013), .CO(N28319), .S(N28318) );
  ad01d0 \add_131_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4793), 
        .B(N4934), .CI(N4928), .CO(N28310), .S(N28309) );
  ad01d0 \add_31_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28157), 
        .B(N27671), .CI(
        \add_31_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_31_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27617)
         );
  ad01d0 \add_31_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28158), 
        .B(N27672), .CI(
        \add_31_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27619), 
        .S(N27618) );
  ad01d0 \add_44_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27869), 
        .B(N27149), .CI(
        \add_44_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27672), 
        .S(N27671) );
  ad01d0 \add_87_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4942), .B(
        N4996), .CI(N4852), .CO(N27869), .S(N27868) );
  ad01d0 \add_43_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27293), 
        .B(N27320), .CI(
        \add_43_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28158), 
        .S(N28157) );
  ad01d0 \add_20_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27716), 
        .B(N27662), .CI(
        \add_20_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_20_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28103)
         );
  ad01d0 \add_20_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27717), 
        .B(N27663), .CI(
        \add_20_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_20_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28104)
         );
  ad01d0 \add_41_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27437), 
        .B(N28400), .CI(
        \add_41_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_41_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27662)
         );
  ad01d0 \add_42_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27284), 
        .B(N27860), .CI(
        \add_42_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28401), 
        .S(N28400) );
  ad01d0 \add_85_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4963), .B(
        N4993), .CI(N4783), .CO(N27860), .S(N27859) );
  ad01d0 \add_53_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27311), 
        .B(N27140), .CI(
        \add_53_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27717), 
        .S(N27716) );
  ad01d0 \add_7_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27536), .B(
        N27545), .CI(\add_7_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_7_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N27500) );
  ad01d0 \add_7_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27537), .B(
        N27546), .CI(\add_7_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_7_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N27501) );
  ad01d0 \add_7_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27538), .B(
        N27547), .CI(\add_7_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_7_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N27502) );
  ad01d0 \add_7_root_add_86_root_add_255_countones_143/U1_4  ( .A(N27539), .B(
        N27548), .CI(\add_7_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(N27504), .S(N27503) );
  ad01d0 \add_16_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28580), 
        .B(N28517), .CI(
        \add_16_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_16_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27545)
         );
  ad01d0 \add_16_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28581), 
        .B(N28518), .CI(
        \add_16_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_16_root_add_86_root_add_255_countones_143/carry[3] ), .S(N27546)
         );
  ad01d0 \add_16_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28582), 
        .B(N28519), .CI(
        \add_16_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N27548), 
        .S(N27547) );
  ad01d0 \add_34_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27779), 
        .B(N27788), .CI(
        \add_34_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_34_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28517)
         );
  ad01d0 \add_34_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27780), 
        .B(N27789), .CI(
        \add_34_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28519), 
        .S(N28518) );
  ad01d0 \add_70_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28337), 
        .B(N27923), .CI(
        \add_70_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27789), 
        .S(N27788) );
  ad01d0 \add_110_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5017), 
        .B(N4876), .CI(N4954), .CO(N27923), .S(N27922) );
  ad01d0 \add_155_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4818), 
        .B(N4821), .CI(N4815), .CO(N28337), .S(N28336) );
  ad01d0 \add_69_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28463), 
        .B(N27203), .CI(
        \add_69_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27780), 
        .S(N27779) );
  ad01d0 \add_108_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4918), 
        .B(N4768), .CI(N4831), .CO(N28463), .S(N28462) );
  ad01d0 \add_33_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27761), 
        .B(N28238), .CI(
        \add_33_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_33_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28580)
         );
  ad01d0 \add_33_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27762), 
        .B(N28239), .CI(
        \add_33_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28582), 
        .S(N28581) );
  ad01d0 \add_78_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27176), 
        .B(N27401), .CI(
        \add_78_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28239), 
        .S(N28238) );
  ad01d0 \add_62_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27275), 
        .B(N28274), .CI(
        \add_62_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27762), 
        .S(N27761) );
  ad01d0 \add_99_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4972), .B(
        N4999), .CI(N4819), .CO(N28274), .S(N28273) );
  ad01d0 \add_14_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27608), 
        .B(N27572), .CI(
        \add_14_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_14_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27536)
         );
  ad01d0 \add_14_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27609), 
        .B(N27573), .CI(
        \add_14_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_14_root_add_86_root_add_255_countones_143/carry[3] ), .S(N27537)
         );
  ad01d0 \add_14_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27610), 
        .B(N27574), .CI(
        \add_14_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N27539), 
        .S(N27538) );
  ad01d0 \add_22_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27698), 
        .B(N28418), .CI(
        \add_22_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_22_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27572)
         );
  ad01d0 \add_22_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27699), 
        .B(N28419), .CI(
        \add_22_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27574), 
        .S(N27573) );
  ad01d0 \add_57_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27878), 
        .B(N27239), .CI(
        \add_57_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28419), 
        .S(N28418) );
  ad01d0 \add_88_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4846), .B(
        N4849), .CI(N4945), .CO(N27878), .S(N27877) );
  ad01d0 \add_48_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27446), 
        .B(N27950), .CI(
        \add_48_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27699), 
        .S(N27698) );
  ad01d0 \add_120_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4856), 
        .B(N4835), .CI(N4988), .CO(N27950), .S(N27949) );
  ad01d0 \add_29_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27743), 
        .B(N27680), .CI(
        \add_29_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_29_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27608)
         );
  ad01d0 \add_29_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27744), 
        .B(N27681), .CI(
        \add_29_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27610), 
        .S(N27609) );
  ad01d0 \add_45_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27995), 
        .B(N27122), .CI(
        \add_45_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27681), 
        .S(N27680) );
  ad01d0 \add_141_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4950), 
        .B(N4881), .CI(N4878), .CO(N27995), .S(N27994) );
  ad01d0 \add_59_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27329), 
        .B(N27383), .CI(
        \add_59_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27744), 
        .S(N27743) );
  ad01d0 \add_6_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27527), .B(
        N28094), .CI(\add_6_root_add_86_root_add_255_countones_143/carry[1] ), 
        .CO(\add_6_root_add_86_root_add_255_countones_143/carry[2] ), .S(
        N27491) );
  ad01d0 \add_6_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27528), .B(
        N28095), .CI(\add_6_root_add_86_root_add_255_countones_143/carry[2] ), 
        .CO(\add_6_root_add_86_root_add_255_countones_143/carry[3] ), .S(
        N27492) );
  ad01d0 \add_6_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27529), .B(
        N28096), .CI(\add_6_root_add_86_root_add_255_countones_143/carry[3] ), 
        .CO(\add_6_root_add_86_root_add_255_countones_143/carry[4] ), .S(
        N27493) );
  ad01d0 \add_6_root_add_86_root_add_255_countones_143/U1_4  ( .A(N27530), .B(
        N28097), .CI(\add_6_root_add_86_root_add_255_countones_143/carry[4] ), 
        .CO(N27495), .S(N27494) );
  ad01d0 \add_15_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27653), 
        .B(N28148), .CI(
        \add_15_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_15_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28094)
         );
  ad01d0 \add_15_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27654), 
        .B(N28149), .CI(
        \add_15_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_15_root_add_86_root_add_255_countones_143/carry[3] ), .S(N28095)
         );
  ad01d0 \add_15_root_add_86_root_add_255_countones_143/U1_3  ( .A(N27655), 
        .B(N28150), .CI(
        \add_15_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N28097), 
        .S(N28096) );
  ad01d0 \add_39_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27824), 
        .B(N28616), .CI(
        \add_39_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_39_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28148)
         );
  ad01d0 \add_39_root_add_86_root_add_255_countones_143/U1_2  ( .A(N27825), 
        .B(N28617), .CI(
        \add_39_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28150), 
        .S(N28149) );
  ad01d0 \add_64_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27887), 
        .B(N27896), .CI(
        \add_64_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28617), 
        .S(N28616) );
  ad01d0 \add_96_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4873), .B(
        N4870), .CI(N4978), .CO(N27896), .S(N27895) );
  ad01d0 \add_93_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4900), .B(
        N4903), .CI(N4975), .CO(N27887), .S(N27886) );
  ad01d0 \add_77_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28004), 
        .B(N27338), .CI(
        \add_77_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N27825), 
        .S(N27824) );
  ad01d0 \add_144_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4866), 
        .B(N4869), .CI(N4863), .CO(N28004), .S(N28003) );
  ad01d0 \add_40_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28445), 
        .B(N28247), .CI(
        \add_40_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_40_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27653)
         );
  ad01d0 \add_40_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28446), 
        .B(N28248), .CI(
        \add_40_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N27655), 
        .S(N27654) );
  ad01d0 \add_83_root_add_86_root_add_255_countones_143/U1_0  ( .A(N27850), 
        .B(N27157), .CI(N4837), .CO(
        \add_83_root_add_86_root_add_255_countones_143/carry[1] ), .S(N28246)
         );
  ad01d0 \add_83_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27851), 
        .B(N27158), .CI(
        \add_83_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28248), 
        .S(N28247) );
  ad01d0 \add_84_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5011), .B(
        N4780), .CI(N4990), .CO(N27851), .S(N27850) );
  ad01d0 \add_82_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28022), 
        .B(N27257), .CI(
        \add_82_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28446), 
        .S(N28445) );
  ad01d0 \add_151_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4833), 
        .B(N4989), .CI(N4938), .CO(N28022), .S(N28021) );
  ad01d0 \add_13_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28130), 
        .B(N28112), .CI(
        \add_13_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_13_root_add_86_root_add_255_countones_143/carry[2] ), .S(N27527)
         );
  ad01d0 \add_13_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28131), 
        .B(N28113), .CI(
        \add_13_root_add_86_root_add_255_countones_143/carry[2] ), .CO(
        \add_13_root_add_86_root_add_255_countones_143/carry[3] ), .S(N27528)
         );
  ad01d0 \add_13_root_add_86_root_add_255_countones_143/U1_3  ( .A(N28132), 
        .B(N28114), .CI(
        \add_13_root_add_86_root_add_255_countones_143/carry[3] ), .CO(N27530), 
        .S(N27529) );
  ad01d0 \add_23_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28409), 
        .B(N28436), .CI(
        \add_23_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_23_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28112)
         );
  ad01d0 \add_23_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28410), 
        .B(N28437), .CI(
        \add_23_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28114), 
        .S(N28113) );
  ad01d0 \add_74_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27194), 
        .B(N28481), .CI(
        \add_74_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28437), 
        .S(N28436) );
  ad01d0 \add_139_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4955), 
        .B(N5018), .CI(N4952), .CO(N28481), .S(N28480) );
  ad01d0 \add_50_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27266), 
        .B(N27959), .CI(
        \add_50_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28410), 
        .S(N28409) );
  ad01d0 \add_125_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4979), 
        .B(N4868), .CI(N4811), .CO(N27959), .S(N27958) );
  ad01d0 \add_30_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28202), 
        .B(N28544), .CI(
        \add_30_root_add_86_root_add_255_countones_143/carry[1] ), .CO(
        \add_30_root_add_86_root_add_255_countones_143/carry[2] ), .S(N28130)
         );
  ad01d0 \add_30_root_add_86_root_add_255_countones_143/U1_2  ( .A(N28203), 
        .B(N28545), .CI(
        \add_30_root_add_86_root_add_255_countones_143/carry[2] ), .CO(N28132), 
        .S(N28131) );
  ad01d0 \add_81_root_add_86_root_add_255_countones_143/U1_1  ( .A(N27905), 
        .B(N28292), .CI(
        \add_81_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28545), 
        .S(N28544) );
  ad01d0 \add_116_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4916), 
        .B(N4853), .CI(N4850), .CO(N28292), .S(N28291) );
  ad01d0 \add_100_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4936), 
        .B(N4879), .CI(N4909), .CO(N27905), .S(N27904) );
  ad01d0 \add_61_root_add_86_root_add_255_countones_143/U1_1  ( .A(N28256), 
        .B(N27392), .CI(
        \add_61_root_add_86_root_add_255_countones_143/carry[1] ), .CO(N28203), 
        .S(N28202) );
  ad01d0 \add_86_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4843), .B(
        N4855), .CI(N4834), .CO(N28256), .S(N28255) );
  ad01d0 \add_168_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4896), 
        .B(N4905), .CI(N4890), .CO(N27482), .S(N27481) );
  ad01d0 \add_167_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4953), 
        .B(N5016), .CI(N4920), .CO(N27473), .S(N27472) );
  ad01d0 \add_165_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5019), 
        .B(N4770), .CI(N4956), .CO(N27464), .S(N27463) );
  ad01d0 \add_164_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4923), 
        .B(N4959), .CI(N4773), .CO(N27455), .S(N27454) );
  ad01d0 \add_161_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4788), 
        .B(N4908), .CI(N4965), .CO(N27446), .S(N27445) );
  ad01d0 \add_160_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4968), 
        .B(N4791), .CI(N4929), .CO(N27437), .S(N27436) );
  ad01d0 \add_158_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4974), 
        .B(N4803), .CI(N4800), .CO(N27428), .S(N27427) );
  ad01d0 \add_157_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4932), 
        .B(N4977), .CI(N4806), .CO(N27419), .S(N27418) );
  ad01d0 \add_153_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4983), 
        .B(N4824), .CI(N4935), .CO(N27410), .S(N27409) );
  ad01d0 \add_152_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4827), 
        .B(N4830), .CI(N4986), .CO(N27401), .S(N27400) );
  ad01d0 \add_150_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4914), 
        .B(N4992), .CI(N4836), .CO(N27392), .S(N27391) );
  ad01d0 \add_149_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4842), 
        .B(N4845), .CI(N4839), .CO(N27383), .S(N27382) );
  ad01d0 \add_146_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4944), 
        .B(N5001), .CI(N4902), .CO(N27374), .S(N27373) );
  ad01d0 \add_145_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4860), 
        .B(N5004), .CI(N4857), .CO(N27365), .S(N27364) );
  ad01d0 \add_143_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4947), 
        .B(N5007), .CI(N4917), .CO(N27356), .S(N27355) );
  ad01d0 \add_142_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5010), 
        .B(N4875), .CI(N4872), .CO(N27347), .S(N27346) );
  ad01d0 \add_137_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4925), 
        .B(N4886), .CI(N4769), .CO(N27338), .S(N27337) );
  ad01d0 \add_136_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4958), 
        .B(N4775), .CI(N4772), .CO(N27329), .S(N27328) );
  ad01d0 \add_134_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4898), 
        .B(N4781), .CI(N4778), .CO(N27320), .S(N27319) );
  ad01d0 \add_133_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4784), 
        .B(N4964), .CI(N5012), .CO(N27311), .S(N27310) );
  ad01d0 \add_130_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4904), 
        .B(N4931), .CI(N4814), .CO(N27302), .S(N27301) );
  ad01d0 \add_129_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4970), 
        .B(N4874), .CI(N4796), .CO(N27293), .S(N27292) );
  ad01d0 \add_127_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4910), 
        .B(N4805), .CI(N4802), .CO(N27284), .S(N27283) );
  ad01d0 \add_126_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4976), 
        .B(N5006), .CI(N4808), .CO(N27275), .S(N27274) );
  ad01d0 \add_122_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4862), 
        .B(N4826), .CI(N4985), .CO(N27266), .S(N27265) );
  ad01d0 \add_121_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4829), 
        .B(N4832), .CI(N4892), .CO(N27257), .S(N27256) );
  ad01d0 \add_119_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5000), 
        .B(N4838), .CI(N4991), .CO(N27248), .S(N27247) );
  ad01d0 \add_118_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4943), 
        .B(N4844), .CI(N4841), .CO(N27239), .S(N27238) );
  ad01d0 \add_115_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5003), 
        .B(N4919), .CI(N4859), .CO(N27230), .S(N27229) );
  ad01d0 \add_114_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4949), 
        .B(N4871), .CI(N4865), .CO(N27221), .S(N27220) );
  ad01d0 \add_112_root_add_86_root_add_255_countones_143/U1_0  ( .A(N5015), 
        .B(N4889), .CI(N4883), .CO(N27212), .S(N27211) );
  ad01d0 \add_111_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4939), 
        .B(N4960), .CI(N4816), .CO(N27203), .S(N27202) );
  ad01d0 \add_105_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4894), 
        .B(N4981), .CI(N4774), .CO(N27194), .S(N27193) );
  ad01d0 \add_104_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4825), 
        .B(N4915), .CI(N5005), .CO(N27185), .S(N27184) );
  ad01d0 \add_102_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4984), 
        .B(N4867), .CI(N4927), .CO(N27176), .S(N27175) );
  ad01d0 \add_101_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4786), 
        .B(N4966), .CI(N4840), .CO(N27167), .S(N27166) );
  ad01d0 \add_98_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4930), .B(
        N4795), .CI(N4807), .CO(N27158), .S(N27157) );
  ad01d0 \add_97_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4798), .B(
        N4813), .CI(N4912), .CO(N27149), .S(N27148) );
  ad01d0 \add_95_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4897), .B(
        N4933), .CI(N4804), .CO(N27140), .S(N27139) );
  ad01d0 \add_94_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4810), .B(
        N4864), .CI(N5008), .CO(N27131), .S(N27130) );
  ad01d0 \add_90_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4792), .B(
        N4858), .CI(N4861), .CO(N27122), .S(N27121) );
  ad01d0 \add_89_root_add_86_root_add_255_countones_143/U1_0  ( .A(N4789), .B(
        N4951), .CI(N4969), .CO(N27113), .S(N27112) );
  dfcrq1 finish_reordering_reg ( .D(n12117), .CP(clk), .CDN(n668), .Q(
        finish_reordering) );
  dfcrq1 new_reference_is_done_reg ( .D(n12189), .CP(clk), .CDN(n584), .Q(
        new_reference_is_done) );
  dfcrq1 \hash_index_reg[1]  ( .D(n2767), .CP(clk), .CDN(n583), .Q(N3877) );
  dfcrq1 \hash_index_reg[2]  ( .D(n12176), .CP(clk), .CDN(n583), .Q(N3878) );
  dfcrq1 distance_ready_reg ( .D(n13793), .CP(clk), .CDN(n586), .Q(
        distance_ready) );
  dfcrq1 finish_flag_reg ( .D(n12203), .CP(clk), .CDN(n592), .Q(finish_flag)
         );
  dfcrq1 reading_current_reg ( .D(n2769), .CP(clk), .CDN(n584), .Q(
        reading_current) );
  dfcrq1 \hash_index_reg[3]  ( .D(n12198), .CP(clk), .CDN(n585), .Q(N3855) );
  dfcrq1 reading_compare_reg ( .D(n12199), .CP(clk), .CDN(n585), .Q(
        reading_compare) );
  dfcrq1 compare_in_progress_reg ( .D(n13794), .CP(clk), .CDN(n584), .Q(
        compare_in_progress) );
  dfcrq1 hashes_ready_reg ( .D(n12200), .CP(clk), .CDN(n586), .Q(hashes_ready)
         );
  dfcrq1 \count_image_reg[8]  ( .D(n12742), .CP(clk), .CDN(n584), .Q(
        count_image[8]) );
  dfcrq1 \compare_image_index_reg[8]  ( .D(n12197), .CP(clk), .CDN(n585), .Q(
        N3182) );
  dfcrq1 \count_image_reg[0]  ( .D(n12741), .CP(clk), .CDN(n584), .Q(
        count_image[0]) );
  dfcrq1 \count_image_reg[1]  ( .D(n12740), .CP(clk), .CDN(n584), .Q(
        count_image[1]) );
  dfcrq1 \images_bus_reg[481]  ( .D(n12772), .CP(clk), .CDN(n591), .Q(
        images_bus[481]) );
  dfcrq1 \compare_image_index_reg[6]  ( .D(n12195), .CP(clk), .CDN(n585), .Q(
        N3180) );
  dfcrq1 \images_bus_reg[225]  ( .D(n13028), .CP(clk), .CDN(n590), .Q(
        images_bus[225]) );
  dfcrq1 \images_bus_reg[449]  ( .D(n12804), .CP(clk), .CDN(n590), .Q(
        images_bus[449]) );
  dfcrq1 \images_bus_reg[483]  ( .D(n12770), .CP(clk), .CDN(n597), .Q(
        images_bus[483]) );
  dfcrq1 \images_bus_reg[236]  ( .D(n13017), .CP(clk), .CDN(n666), .Q(
        images_bus[236]) );
  dfcrq1 \images_bus_reg[485]  ( .D(n12768), .CP(clk), .CDN(n579), .Q(
        images_bus[485]) );
  dfcrq1 \images_bus_reg[193]  ( .D(n13060), .CP(clk), .CDN(n590), .Q(
        images_bus[193]) );
  dfcrq1 \images_bus_reg[451]  ( .D(n12802), .CP(clk), .CDN(n597), .Q(
        images_bus[451]) );
  dfcrq1 \images_bus_reg[246]  ( .D(n13007), .CP(clk), .CDN(n557), .Q(
        images_bus[246]) );
  dfcrq1 \images_bus_reg[196]  ( .D(n13057), .CP(clk), .CDN(n573), .Q(
        images_bus[196]) );
  dfcrq1 \images_bus_reg[161]  ( .D(n13092), .CP(clk), .CDN(n590), .Q(
        images_bus[161]) );
  dfcrq1 \images_bus_reg[457]  ( .D(n12796), .CP(clk), .CDN(n592), .Q(
        images_bus[457]) );
  dfcrq1 \images_bus_reg[505]  ( .D(n12748), .CP(clk), .CDN(n595), .Q(
        images_bus[505]) );
  dfcrq1 \images_bus_reg[241]  ( .D(n13012), .CP(clk), .CDN(n593), .Q(
        images_bus[241]) );
  dfcrq1 \images_bus_reg[417]  ( .D(n12836), .CP(clk), .CDN(n590), .Q(
        images_bus[417]) );
  dfcrq1 \images_bus_reg[456]  ( .D(n12797), .CP(clk), .CDN(n564), .Q(
        images_bus[456]) );
  dfcrq1 \images_bus_reg[252]  ( .D(n13001), .CP(clk), .CDN(n553), .Q(
        images_bus[252]) );
  dfcrq1 \images_bus_reg[230]  ( .D(n13023), .CP(clk), .CDN(n554), .Q(
        images_bus[230]) );
  dfcrq1 \images_bus_reg[488]  ( .D(n12765), .CP(clk), .CDN(n564), .Q(
        images_bus[488]) );
  dfcrq1 \images_bus_reg[238]  ( .D(n13015), .CP(clk), .CDN(n555), .Q(
        images_bus[238]) );
  dfcrq1 \images_bus_reg[243]  ( .D(n13010), .CP(clk), .CDN(n575), .Q(
        images_bus[243]) );
  dfcrq1 \images_bus_reg[453]  ( .D(n12800), .CP(clk), .CDN(n578), .Q(
        images_bus[453]) );
  dfcrq1 \images_bus_reg[480]  ( .D(n12773), .CP(clk), .CDN(n563), .Q(
        images_bus[480]) );
  dfcrq1 \images_bus_reg[224]  ( .D(n13029), .CP(clk), .CDN(n562), .Q(
        images_bus[224]) );
  dfcrq1 \images_bus_reg[229]  ( .D(n13024), .CP(clk), .CDN(n578), .Q(
        images_bus[229]) );
  dfcrq1 \images_bus_reg[244]  ( .D(n13009), .CP(clk), .CDN(n551), .Q(
        images_bus[244]) );
  dfcrq1 \images_bus_reg[385]  ( .D(n12868), .CP(clk), .CDN(n590), .Q(
        images_bus[385]) );
  dfcrq1 \images_bus_reg[454]  ( .D(n12799), .CP(clk), .CDN(n554), .Q(
        images_bus[454]) );
  dfcrq1 \images_bus_reg[172]  ( .D(n13081), .CP(clk), .CDN(n704), .Q(
        images_bus[172]) );
  dfcrq1 \images_bus_reg[201]  ( .D(n13052), .CP(clk), .CDN(n591), .Q(
        images_bus[201]) );
  dfcrq1 \images_bus_reg[203]  ( .D(n13050), .CP(clk), .CDN(n597), .Q(
        images_bus[203]) );
  dfcrq1 \images_bus_reg[486]  ( .D(n12767), .CP(clk), .CDN(n555), .Q(
        images_bus[486]) );
  dfcrq1 \images_bus_reg[487]  ( .D(n12766), .CP(clk), .CDN(n586), .Q(
        images_bus[487]) );
  dfcrq1 \images_bus_reg[387]  ( .D(n12866), .CP(clk), .CDN(n596), .Q(
        images_bus[387]) );
  dfcrq1 \images_bus_reg[198]  ( .D(n13055), .CP(clk), .CDN(n554), .Q(
        images_bus[198]) );
  dfcrq1 \images_bus_reg[398]  ( .D(n12855), .CP(clk), .CDN(n556), .Q(
        images_bus[398]) );
  dfcrq1 \images_bus_reg[177]  ( .D(n13076), .CP(clk), .CDN(n593), .Q(
        images_bus[177]) );
  dfcrq1 \images_bus_reg[499]  ( .D(n12754), .CP(clk), .CDN(n576), .Q(
        images_bus[499]) );
  dfcrq1 \images_bus_reg[460]  ( .D(n12793), .CP(clk), .CDN(n551), .Q(
        images_bus[460]) );
  dfcrq1 \count_image_reg[2]  ( .D(n12739), .CP(clk), .CDN(n584), .Q(
        count_image[2]) );
  dfcrq1 \images_bus_reg[145]  ( .D(n13108), .CP(clk), .CDN(n592), .Q(
        images_bus[145]) );
  dfcrq1 \images_bus_reg[491]  ( .D(n12762), .CP(clk), .CDN(n574), .Q(
        images_bus[491]) );
  dfcrq1 \images_bus_reg[165]  ( .D(n13088), .CP(clk), .CDN(n578), .Q(
        images_bus[165]) );
  dfcrq1 \images_bus_reg[459]  ( .D(n12794), .CP(clk), .CDN(n574), .Q(
        images_bus[459]) );
  dfcrq1 \images_bus_reg[192]  ( .D(n13061), .CP(clk), .CDN(n562), .Q(
        images_bus[192]) );
  dfcrq1 \images_bus_reg[212]  ( .D(n13041), .CP(clk), .CDN(n551), .Q(
        images_bus[212]) );
  dfcrq1 \images_bus_reg[233]  ( .D(n13020), .CP(clk), .CDN(n591), .Q(
        images_bus[233]) );
  dfcrq1 \images_bus_reg[419]  ( .D(n12834), .CP(clk), .CDN(n596), .Q(
        images_bus[419]) );
  dfcrq1 \images_bus_reg[436]  ( .D(n12817), .CP(clk), .CDN(n552), .Q(
        images_bus[436]) );
  dfcrq1 \images_bus_reg[493]  ( .D(n12760), .CP(clk), .CDN(n580), .Q(
        images_bus[493]) );
  dfcrq1 \images_bus_reg[500]  ( .D(n12753), .CP(clk), .CDN(n552), .Q(
        images_bus[500]) );
  dfcrq1 \images_bus_reg[450]  ( .D(n12803), .CP(clk), .CDN(n569), .Q(
        images_bus[450]) );
  dfcrq1 \images_bus_reg[425]  ( .D(n12828), .CP(clk), .CDN(n592), .Q(
        images_bus[425]) );
  dfcrq1 \images_bus_reg[227]  ( .D(n13026), .CP(clk), .CDN(n596), .Q(
        images_bus[227]) );
  dfcrq1 \images_bus_reg[506]  ( .D(n12747), .CP(clk), .CDN(n572), .Q(
        images_bus[506]) );
  dfcrq1 \images_bus_reg[231]  ( .D(n13022), .CP(clk), .CDN(n561), .Q(
        images_bus[231]) );
  dfcrq1 \images_bus_reg[195]  ( .D(n13058), .CP(clk), .CDN(n596), .Q(
        images_bus[195]) );
  dfcrq1 \images_bus_reg[497]  ( .D(n12756), .CP(clk), .CDN(n594), .Q(
        images_bus[497]) );
  dfcrq1 \images_bus_reg[142]  ( .D(n13111), .CP(clk), .CDN(n555), .Q(
        images_bus[142]) );
  dfcrq1 \images_bus_reg[467]  ( .D(n12786), .CP(clk), .CDN(n576), .Q(
        images_bus[467]) );
  dfcrq1 \images_bus_reg[509]  ( .D(n12744), .CP(clk), .CDN(n583), .Q(
        images_bus[509]) );
  dfcrq1 \images_bus_reg[245]  ( .D(n13008), .CP(clk), .CDN(n581), .Q(
        images_bus[245]) );
  dfcrq1 \images_bus_reg[137]  ( .D(n13116), .CP(clk), .CDN(n591), .Q(
        images_bus[137]) );
  dfcrq1 \images_bus_reg[36]  ( .D(n13217), .CP(clk), .CDN(n573), .Q(
        images_bus[36]) );
  dfcrq1 \images_bus_reg[217]  ( .D(n13036), .CP(clk), .CDN(n594), .Q(
        images_bus[217]) );
  dfcrq1 \images_bus_reg[97]  ( .D(n13156), .CP(clk), .CDN(n589), .Q(
        images_bus[97]) );
  dfcrq1 \images_bus_reg[393]  ( .D(n12860), .CP(clk), .CDN(n592), .Q(
        images_bus[393]) );
  dfcrq1 \images_bus_reg[321]  ( .D(n12932), .CP(clk), .CDN(n590), .Q(
        images_bus[321]) );
  dfcrq1 \images_bus_reg[422]  ( .D(n12831), .CP(clk), .CDN(n554), .Q(
        images_bus[422]) );
  dfcrq1 \images_bus_reg[473]  ( .D(n12780), .CP(clk), .CDN(n595), .Q(
        images_bus[473]) );
  dfcrq1 \images_bus_reg[490]  ( .D(n12763), .CP(clk), .CDN(n570), .Q(
        images_bus[490]) );
  dfcrq1 \images_bus_reg[209]  ( .D(n13044), .CP(clk), .CDN(n593), .Q(
        images_bus[209]) );
  dfcrq1 \images_bus_reg[353]  ( .D(n12900), .CP(clk), .CDN(n590), .Q(
        images_bus[353]) );
  dfcrq1 \images_bus_reg[100]  ( .D(n13153), .CP(clk), .CDN(n573), .Q(
        images_bus[100]) );
  dfcrq1 \images_bus_reg[129]  ( .D(n13124), .CP(clk), .CDN(n589), .Q(
        images_bus[129]) );
  dfcrq1 \images_bus_reg[134]  ( .D(n13119), .CP(clk), .CDN(n554), .Q(
        images_bus[134]) );
  dfcrq1 \images_bus_reg[455]  ( .D(n12798), .CP(clk), .CDN(n562), .Q(
        images_bus[455]) );
  dfcrq1 \images_bus_reg[215]  ( .D(n13038), .CP(clk), .CDN(n588), .Q(
        images_bus[215]) );
  dfcrq1 \images_bus_reg[424]  ( .D(n12829), .CP(clk), .CDN(n564), .Q(
        images_bus[424]) );
  dfcrq1 \images_bus_reg[164]  ( .D(n13089), .CP(clk), .CDN(n573), .Q(
        images_bus[164]) );
  dfcrq1 \images_bus_reg[498]  ( .D(n12755), .CP(clk), .CDN(n571), .Q(
        images_bus[498]) );
  dfcrq1 \images_bus_reg[240]  ( .D(n13013), .CP(clk), .CDN(n565), .Q(
        images_bus[240]) );
  dfcrq1 \images_bus_reg[128]  ( .D(n13125), .CP(clk), .CDN(n562), .Q(
        images_bus[128]) );
  dfcrq1 \images_bus_reg[200]  ( .D(n13053), .CP(clk), .CDN(n564), .Q(
        images_bus[200]) );
  dfcrq1 \images_bus_reg[234]  ( .D(n13019), .CP(clk), .CDN(n569), .Q(
        images_bus[234]) );
  dfcrq1 \images_bus_reg[484]  ( .D(n12769), .CP(clk), .CDN(n573), .Q(
        images_bus[484]) );
  dfcrq1 \images_bus_reg[471]  ( .D(n12782), .CP(clk), .CDN(n589), .Q(
        images_bus[471]) );
  dfcrq1 \images_bus_reg[162]  ( .D(n13091), .CP(clk), .CDN(n568), .Q(
        images_bus[162]) );
  dfcrq1 \images_bus_reg[160]  ( .D(n13093), .CP(clk), .CDN(n562), .Q(
        images_bus[160]) );
  dfcrq1 \images_bus_reg[433]  ( .D(n12820), .CP(clk), .CDN(n593), .Q(
        images_bus[433]) );
  dfcrq1 \images_bus_reg[435]  ( .D(n12818), .CP(clk), .CDN(n575), .Q(
        images_bus[435]) );
  dfcrq1 \images_bus_reg[492]  ( .D(n12761), .CP(clk), .CDN(n551), .Q(
        images_bus[492]) );
  dfcrq1 \images_bus_reg[33]  ( .D(n13220), .CP(clk), .CDN(n589), .Q(
        images_bus[33]) );
  dfcrq1 \images_bus_reg[475]  ( .D(n12778), .CP(clk), .CDN(n577), .Q(
        images_bus[475]) );
  dfcrq1 \images_bus_reg[99]  ( .D(n13154), .CP(clk), .CDN(n595), .Q(
        images_bus[99]) );
  dfcrq1 \images_bus_reg[507]  ( .D(n12746), .CP(clk), .CDN(n577), .Q(
        images_bus[507]) );
  dfcrq1 \images_bus_reg[461]  ( .D(n12792), .CP(clk), .CDN(n580), .Q(
        images_bus[461]) );
  dfcrq1 \images_bus_reg[131]  ( .D(n13122), .CP(clk), .CDN(n596), .Q(
        images_bus[131]) );
  dfcrq1 \images_bus_reg[502]  ( .D(n12751), .CP(clk), .CDN(n557), .Q(
        images_bus[502]) );
  dfcrq1 \images_bus_reg[401]  ( .D(n12852), .CP(clk), .CDN(n593), .Q(
        images_bus[401]) );
  dfcrq1 \images_bus_reg[211]  ( .D(n13042), .CP(clk), .CDN(n575), .Q(
        images_bus[211]) );
  dfcrq1 \images_bus_reg[68]  ( .D(n13185), .CP(clk), .CDN(n573), .Q(
        images_bus[68]) );
  dfcrq1 \images_bus_reg[503]  ( .D(n12750), .CP(clk), .CDN(n589), .Q(
        images_bus[503]) );
  dfcrq1 \images_bus_reg[465]  ( .D(n12788), .CP(clk), .CDN(n593), .Q(
        images_bus[465]) );
  dfcrq1 \images_bus_reg[171]  ( .D(n13082), .CP(clk), .CDN(n597), .Q(
        images_bus[171]) );
  dfcrq1 \images_bus_reg[389]  ( .D(n12864), .CP(clk), .CDN(n578), .Q(
        images_bus[389]) );
  dfcrq1 \images_bus_reg[188]  ( .D(n13065), .CP(clk), .CDN(n552), .Q(
        images_bus[188]) );
  dfcrq1 \images_bus_reg[437]  ( .D(n12816), .CP(clk), .CDN(n581), .Q(
        images_bus[437]) );
  dfcrq1 \images_bus_reg[242]  ( .D(n13011), .CP(clk), .CDN(n570), .Q(
        images_bus[242]) );
  dfcrq1 \images_bus_reg[199]  ( .D(n13054), .CP(clk), .CDN(n561), .Q(
        images_bus[199]) );
  dfcrq1 \images_bus_reg[390]  ( .D(n12863), .CP(clk), .CDN(n554), .Q(
        images_bus[390]) );
  dfcrq1 \images_bus_reg[251]  ( .D(n13002), .CP(clk), .CDN(n576), .Q(
        images_bus[251]) );
  dfcrq1 \images_bus_reg[3]  ( .D(n13250), .CP(clk), .CDN(n595), .Q(
        images_bus[3]) );
  dfcrq1 \images_bus_reg[65]  ( .D(n13188), .CP(clk), .CDN(n589), .Q(
        images_bus[65]) );
  dfcrq1 \images_bus_reg[214]  ( .D(n13039), .CP(clk), .CDN(n557), .Q(
        images_bus[214]) );
  dfcrq1 \images_bus_reg[253]  ( .D(n13000), .CP(clk), .CDN(n582), .Q(
        images_bus[253]) );
  dfcrq1 \images_bus_reg[249]  ( .D(n13004), .CP(clk), .CDN(n594), .Q(
        images_bus[249]) );
  dfcrq1 \images_bus_reg[169]  ( .D(n13084), .CP(clk), .CDN(n591), .Q(
        images_bus[169]) );
  dfcrq1 \images_bus_reg[213]  ( .D(n13040), .CP(clk), .CDN(n581), .Q(
        images_bus[213]) );
  dfcrq1 \images_bus_reg[429]  ( .D(n12824), .CP(clk), .CDN(n580), .Q(
        images_bus[429]) );
  dfcrq1 \images_bus_reg[173]  ( .D(n13080), .CP(clk), .CDN(n579), .Q(
        images_bus[173]) );
  dfcrq1 \images_bus_reg[163]  ( .D(n13090), .CP(clk), .CDN(n596), .Q(
        images_bus[163]) );
  dfcrq1 \images_bus_reg[472]  ( .D(n12781), .CP(clk), .CDN(n567), .Q(
        images_bus[472]) );
  dfcrq1 \images_bus_reg[181]  ( .D(n13072), .CP(clk), .CDN(n581), .Q(
        images_bus[181]) );
  dfcrq1 \images_bus_reg[423]  ( .D(n12830), .CP(clk), .CDN(n561), .Q(
        images_bus[423]) );
  dfcrq1 \images_bus_reg[426]  ( .D(n12827), .CP(clk), .CDN(n570), .Q(
        images_bus[426]) );
  dfcrq1 \count_image_reg[6]  ( .D(n12735), .CP(clk), .CDN(n584), .Q(
        count_image[6]) );
  dfcrq1 \images_bus_reg[237]  ( .D(n13016), .CP(clk), .CDN(n579), .Q(
        images_bus[237]) );
  dfcrq1 \images_bus_reg[395]  ( .D(n12858), .CP(clk), .CDN(n574), .Q(
        images_bus[395]) );
  dfcrq1 \images_bus_reg[35]  ( .D(n13218), .CP(clk), .CDN(n595), .Q(
        images_bus[35]) );
  dfcrq1 \images_bus_reg[392]  ( .D(n12861), .CP(clk), .CDN(n564), .Q(
        images_bus[392]) );
  dfcrq1 \images_bus_reg[430]  ( .D(n12823), .CP(clk), .CDN(n556), .Q(
        images_bus[430]) );
  dfcrq1 \images_bus_reg[220]  ( .D(n13033), .CP(clk), .CDN(n553), .Q(
        images_bus[220]) );
  dfcrq1 \images_bus_reg[166]  ( .D(n13087), .CP(clk), .CDN(n554), .Q(
        images_bus[166]) );
  dfcrq1 \images_bus_reg[194]  ( .D(n13059), .CP(clk), .CDN(n568), .Q(
        images_bus[194]) );
  dfcrq1 \images_bus_reg[235]  ( .D(n13018), .CP(clk), .CDN(n597), .Q(
        images_bus[235]) );
  dfcrq1 \images_bus_reg[384]  ( .D(n12869), .CP(clk), .CDN(n563), .Q(
        images_bus[384]) );
  dfcrq1 \images_bus_reg[141]  ( .D(n13112), .CP(clk), .CDN(n579), .Q(
        images_bus[141]) );
  dfcrq1 \images_bus_reg[179]  ( .D(n13074), .CP(clk), .CDN(n575), .Q(
        images_bus[179]) );
  dfcrq1 \images_bus_reg[396]  ( .D(n12857), .CP(clk), .CDN(n551), .Q(
        images_bus[396]) );
  dfcrq1 \images_bus_reg[444]  ( .D(n12809), .CP(clk), .CDN(n553), .Q(
        images_bus[444]) );
  dfcrq1 \images_bus_reg[250]  ( .D(n13003), .CP(clk), .CDN(n572), .Q(
        images_bus[250]) );
  dfcrq1 \images_bus_reg[176]  ( .D(n13077), .CP(clk), .CDN(n565), .Q(
        images_bus[176]) );
  dfcrq1 \images_bus_reg[147]  ( .D(n13106), .CP(clk), .CDN(n575), .Q(
        images_bus[147]) );
  dfcrq1 \images_bus_reg[466]  ( .D(n12787), .CP(clk), .CDN(n571), .Q(
        images_bus[466]) );
  dfcrq1 \images_bus_reg[248]  ( .D(n13005), .CP(clk), .CDN(n567), .Q(
        images_bus[248]) );
  dfcrq1 \images_bus_reg[219]  ( .D(n13034), .CP(clk), .CDN(n576), .Q(
        images_bus[219]) );
  dfcrq1 \images_bus_reg[102]  ( .D(n13151), .CP(clk), .CDN(n553), .Q(
        images_bus[102]) );
  dfcrq1 \images_bus_reg[208]  ( .D(n13045), .CP(clk), .CDN(n565), .Q(
        images_bus[208]) );
  dfcrq1 \images_bus_reg[494]  ( .D(n12759), .CP(clk), .CDN(n556), .Q(
        images_bus[494]) );
  dfcrq1 \images_bus_reg[477]  ( .D(n12776), .CP(clk), .CDN(n583), .Q(
        images_bus[477]) );
  dfcrq1 \images_bus_reg[185]  ( .D(n13068), .CP(clk), .CDN(n594), .Q(
        images_bus[185]) );
  dfcrq1 \images_bus_reg[427]  ( .D(n12826), .CP(clk), .CDN(n574), .Q(
        images_bus[427]) );
  dfcrq1 \images_bus_reg[496]  ( .D(n12757), .CP(clk), .CDN(n566), .Q(
        images_bus[496]) );
  dfcrq1 \images_bus_reg[365]  ( .D(n12888), .CP(clk), .CDN(n580), .Q(
        images_bus[365]) );
  dfcrq1 \images_bus_reg[52]  ( .D(n13201), .CP(clk), .CDN(n551), .Q(
        images_bus[52]) );
  dfcrq1 \images_bus_reg[124]  ( .D(n13129), .CP(clk), .CDN(n552), .Q(
        images_bus[124]) );
  dfcrq1 \images_bus_reg[355]  ( .D(n12898), .CP(clk), .CDN(n596), .Q(
        images_bus[355]) );
  dfcrq1 \images_bus_reg[5]  ( .D(n13248), .CP(clk), .CDN(n577), .Q(
        images_bus[5]) );
  dfcrq1 \images_bus_reg[216]  ( .D(n13037), .CP(clk), .CDN(n567), .Q(
        images_bus[216]) );
  dfcrq1 \images_bus_reg[418]  ( .D(n12835), .CP(clk), .CDN(n569), .Q(
        images_bus[418]) );
  dfcrq1 \images_bus_reg[149]  ( .D(n13104), .CP(clk), .CDN(n581), .Q(
        images_bus[149]) );
  dfcrq1 \images_bus_reg[133]  ( .D(n13120), .CP(clk), .CDN(n578), .Q(
        images_bus[133]) );
  dfcrq1 \images_bus_reg[1]  ( .D(n13252), .CP(clk), .CDN(n589), .Q(
        images_bus[1]) );
  dfcrq1 \images_bus_reg[113]  ( .D(n13140), .CP(clk), .CDN(n592), .Q(
        images_bus[113]) );
  dfcrq1 \images_bus_reg[210]  ( .D(n13043), .CP(clk), .CDN(n570), .Q(
        images_bus[210]) );
  dfcrq1 \images_bus_reg[369]  ( .D(n12884), .CP(clk), .CDN(n593), .Q(
        images_bus[369]) );
  dfcrq1 \images_bus_reg[221]  ( .D(n13032), .CP(clk), .CDN(n582), .Q(
        images_bus[221]) );
  dfcrq1 \images_bus_reg[495]  ( .D(n12758), .CP(clk), .CDN(n587), .Q(
        images_bus[495]) );
  dfcrq1 \images_bus_reg[130]  ( .D(n13123), .CP(clk), .CDN(n568), .Q(
        images_bus[130]) );
  dfcrq1 \images_bus_reg[254]  ( .D(n12999), .CP(clk), .CDN(n558), .Q(
        images_bus[254]) );
  dfcrq1 \images_bus_reg[205]  ( .D(n13048), .CP(clk), .CDN(n579), .Q(
        images_bus[205]) );
  dfcrq1 \images_bus_reg[255]  ( .D(n12998), .CP(clk), .CDN(n559), .Q(
        images_bus[255]) );
  dfcrq1 \images_bus_reg[135]  ( .D(n13118), .CP(clk), .CDN(n561), .Q(
        images_bus[135]) );
  dfcrq1 \images_bus_reg[421]  ( .D(n12832), .CP(clk), .CDN(n578), .Q(
        images_bus[421]) );
  dfcrq1 \images_bus_reg[443]  ( .D(n12810), .CP(clk), .CDN(n577), .Q(
        images_bus[443]) );
  dfcrq1 \images_bus_reg[81]  ( .D(n13172), .CP(clk), .CDN(n592), .Q(
        images_bus[81]) );
  dfcrq1 \images_bus_reg[372]  ( .D(n12881), .CP(clk), .CDN(n552), .Q(
        images_bus[372]) );
  dfcrq1 \images_bus_reg[292]  ( .D(n12961), .CP(clk), .CDN(n573), .Q(
        images_bus[292]) );
  dfcrq1 \images_bus_reg[132]  ( .D(n13121), .CP(clk), .CDN(n573), .Q(
        images_bus[132]) );
  dfcrq1 \images_bus_reg[411]  ( .D(n12842), .CP(clk), .CDN(n577), .Q(
        images_bus[411]) );
  dfcrq1 \images_bus_reg[448]  ( .D(n12805), .CP(clk), .CDN(n563), .Q(
        images_bus[448]) );
  dfcrq1 \images_bus_reg[405]  ( .D(n12848), .CP(clk), .CDN(n581), .Q(
        images_bus[405]) );
  dfcrq1 \images_bus_reg[414]  ( .D(n12839), .CP(clk), .CDN(n559), .Q(
        images_bus[414]) );
  dfcrq1 \images_bus_reg[153]  ( .D(n13100), .CP(clk), .CDN(n594), .Q(
        images_bus[153]) );
  dfcrq1 \images_bus_reg[431]  ( .D(n12822), .CP(clk), .CDN(n587), .Q(
        images_bus[431]) );
  dfcrq1 \images_bus_reg[357]  ( .D(n12896), .CP(clk), .CDN(n578), .Q(
        images_bus[357]) );
  dfcrq1 \images_bus_reg[110]  ( .D(n13143), .CP(clk), .CDN(n555), .Q(
        images_bus[110]) );
  dfcrq1 \images_bus_reg[504]  ( .D(n12749), .CP(clk), .CDN(n568), .Q(
        images_bus[504]) );
  dfcrq1 \images_bus_reg[144]  ( .D(n13109), .CP(clk), .CDN(n565), .Q(
        images_bus[144]) );
  dfcrq1 \images_bus_reg[170]  ( .D(n13083), .CP(clk), .CDN(n569), .Q(
        images_bus[170]) );
  dfcrq1 \images_bus_reg[440]  ( .D(n12813), .CP(clk), .CDN(n567), .Q(
        images_bus[440]) );
  dfcrq1 \images_bus_reg[325]  ( .D(n12928), .CP(clk), .CDN(n578), .Q(
        images_bus[325]) );
  dfcrq1 \images_bus_reg[469]  ( .D(n12784), .CP(clk), .CDN(n582), .Q(
        images_bus[469]) );
  dfcrq1 \images_bus_reg[155]  ( .D(n13098), .CP(clk), .CDN(n576), .Q(
        images_bus[155]) );
  dfcrq1 \images_bus_reg[394]  ( .D(n12859), .CP(clk), .CDN(n570), .Q(
        images_bus[394]) );
  dfcrq1 \images_bus_reg[80]  ( .D(n13173), .CP(clk), .CDN(n565), .Q(
        images_bus[80]) );
  dfcrq1 \images_bus_reg[151]  ( .D(n13102), .CP(clk), .CDN(n588), .Q(
        images_bus[151]) );
  dfcrq1 \images_bus_reg[4]  ( .D(n13249), .CP(clk), .CDN(n572), .Q(
        images_bus[4]) );
  dfcrq1 \images_bus_reg[289]  ( .D(n12964), .CP(clk), .CDN(n590), .Q(
        images_bus[289]) );
  dfcrq1 \images_bus_reg[320]  ( .D(n12933), .CP(clk), .CDN(n562), .Q(
        images_bus[320]) );
  dfcrq1 \images_bus_reg[49]  ( .D(n13204), .CP(clk), .CDN(n592), .Q(
        images_bus[49]) );
  dfcrq1 \images_bus_reg[464]  ( .D(n12789), .CP(clk), .CDN(n566), .Q(
        images_bus[464]) );
  dfcrq1 \images_bus_reg[73]  ( .D(n13180), .CP(clk), .CDN(n591), .Q(
        images_bus[73]) );
  dfcrq1 \images_bus_reg[445]  ( .D(n12808), .CP(clk), .CDN(n583), .Q(
        images_bus[445]) );
  dfcrq1 \images_bus_reg[107]  ( .D(n13146), .CP(clk), .CDN(n597), .Q(
        images_bus[107]) );
  dfcrq1 \images_bus_reg[108]  ( .D(n13145), .CP(clk), .CDN(n549), .Q(
        images_bus[108]) );
  dfcrq1 \images_bus_reg[67]  ( .D(n13186), .CP(clk), .CDN(n595), .Q(
        images_bus[67]) );
  dfcrq1 \images_bus_reg[43]  ( .D(n13210), .CP(clk), .CDN(n597), .Q(
        images_bus[43]) );
  dfcrq1 \images_bus_reg[178]  ( .D(n13075), .CP(clk), .CDN(n570), .Q(
        images_bus[178]) );
  dfcrq1 \images_bus_reg[118]  ( .D(n13135), .CP(clk), .CDN(n556), .Q(
        images_bus[118]) );
  dfcrq1 \images_bus_reg[39]  ( .D(n13214), .CP(clk), .CDN(n560), .Q(
        images_bus[39]) );
  dfcrq1 \images_bus_reg[75]  ( .D(n13178), .CP(clk), .CDN(n597), .Q(
        images_bus[75]) );
  dfcrq1 \images_bus_reg[140]  ( .D(n13113), .CP(clk), .CDN(n546), .Q(
        images_bus[140]) );
  dfcrq1 \images_bus_reg[112]  ( .D(n13141), .CP(clk), .CDN(n565), .Q(
        images_bus[112]) );
  dfcrq1 \images_bus_reg[261]  ( .D(n12992), .CP(clk), .CDN(n578), .Q(
        images_bus[261]) );
  dfcrq1 \images_bus_reg[189]  ( .D(n13064), .CP(clk), .CDN(n582), .Q(
        images_bus[189]) );
  dfcrq1 \images_bus_reg[167]  ( .D(n13086), .CP(clk), .CDN(n561), .Q(
        images_bus[167]) );
  dfcrq1 \images_bus_reg[413]  ( .D(n12840), .CP(clk), .CDN(n583), .Q(
        images_bus[413]) );
  dfcrq1 \images_bus_reg[150]  ( .D(n13103), .CP(clk), .CDN(n556), .Q(
        images_bus[150]) );
  dfcrq1 \images_bus_reg[98]  ( .D(n13155), .CP(clk), .CDN(n568), .Q(
        images_bus[98]) );
  dfcrq1 \images_bus_reg[96]  ( .D(n13157), .CP(clk), .CDN(n562), .Q(
        images_bus[96]) );
  dfcrq1 \images_bus_reg[260]  ( .D(n12993), .CP(clk), .CDN(n573), .Q(
        images_bus[260]) );
  dfcrq1 \images_bus_reg[186]  ( .D(n13067), .CP(clk), .CDN(n572), .Q(
        images_bus[186]) );
  dfcrq1 \images_bus_reg[183]  ( .D(n13070), .CP(clk), .CDN(n588), .Q(
        images_bus[183]) );
  dfcrq1 \images_bus_reg[83]  ( .D(n13170), .CP(clk), .CDN(n574), .Q(
        images_bus[83]) );
  dfcrq1 \images_bus_reg[191]  ( .D(n13062), .CP(clk), .CDN(n559), .Q(
        images_bus[191]) );
  dfcrq1 \images_bus_reg[442]  ( .D(n12811), .CP(clk), .CDN(n572), .Q(
        images_bus[442]) );
  dfcrq1 \images_bus_reg[329]  ( .D(n12924), .CP(clk), .CDN(n592), .Q(
        images_bus[329]) );
  dfcrq1 \images_bus_reg[78]  ( .D(n13175), .CP(clk), .CDN(n555), .Q(
        images_bus[78]) );
  dfcrq1 \images_bus_reg[101]  ( .D(n13152), .CP(clk), .CDN(n577), .Q(
        images_bus[101]) );
  dfcrq1 \images_bus_reg[158]  ( .D(n13095), .CP(clk), .CDN(n558), .Q(
        images_bus[158]) );
  dfcrq1 \images_bus_reg[377]  ( .D(n12876), .CP(clk), .CDN(n595), .Q(
        images_bus[377]) );
  dfcrq1 \images_bus_reg[247]  ( .D(n13006), .CP(clk), .CDN(n588), .Q(
        images_bus[247]) );
  dfcrq1 \images_bus_reg[204]  ( .D(n13049), .CP(clk), .CDN(n707), .Q(
        images_bus[204]) );
  dfcrq1 \images_bus_reg[109]  ( .D(n13144), .CP(clk), .CDN(n579), .Q(
        images_bus[109]) );
  dfcrq1 \images_bus_reg[409]  ( .D(n12844), .CP(clk), .CDN(n595), .Q(
        images_bus[409]) );
  dfcrq1 \images_bus_reg[72]  ( .D(n13181), .CP(clk), .CDN(n563), .Q(
        images_bus[72]) );
  dfcrq1 \images_bus_reg[37]  ( .D(n13216), .CP(clk), .CDN(n577), .Q(
        images_bus[37]) );
  dfcrq1 \images_bus_reg[115]  ( .D(n13138), .CP(clk), .CDN(n574), .Q(
        images_bus[115]) );
  dfcrq1 \images_bus_reg[156]  ( .D(n13097), .CP(clk), .CDN(n552), .Q(
        images_bus[156]) );
  dfcrq1 \images_bus_reg[38]  ( .D(n13215), .CP(clk), .CDN(n553), .Q(
        images_bus[38]) );
  dfcrq1 \images_bus_reg[447]  ( .D(n12806), .CP(clk), .CDN(n560), .Q(
        images_bus[447]) );
  dfcrq1 \images_bus_reg[84]  ( .D(n13169), .CP(clk), .CDN(n551), .Q(
        images_bus[84]) );
  dfcrq1 \images_bus_reg[434]  ( .D(n12819), .CP(clk), .CDN(n571), .Q(
        images_bus[434]) );
  dfcrq1 \images_bus_reg[416]  ( .D(n12837), .CP(clk), .CDN(n563), .Q(
        images_bus[416]) );
  dfcrq1 \images_bus_reg[474]  ( .D(n12779), .CP(clk), .CDN(n572), .Q(
        images_bus[474]) );
  dfcrq1 \images_bus_reg[352]  ( .D(n12901), .CP(clk), .CDN(n563), .Q(
        images_bus[352]) );
  dfcrq1 \images_bus_reg[403]  ( .D(n12850), .CP(clk), .CDN(n575), .Q(
        images_bus[403]) );
  dfcrq1 \images_bus_reg[391]  ( .D(n12862), .CP(clk), .CDN(n561), .Q(
        images_bus[391]) );
  dfcrq1 \images_bus_reg[337]  ( .D(n12916), .CP(clk), .CDN(n593), .Q(
        images_bus[337]) );
  dfcrq1 \images_bus_reg[408]  ( .D(n12845), .CP(clk), .CDN(n567), .Q(
        images_bus[408]) );
  dfcrq1 \images_bus_reg[406]  ( .D(n12847), .CP(clk), .CDN(n557), .Q(
        images_bus[406]) );
  dfcrq1 \images_bus_reg[463]  ( .D(n12790), .CP(clk), .CDN(n587), .Q(
        images_bus[463]) );
  dfcrq1 \images_bus_reg[111]  ( .D(n13142), .CP(clk), .CDN(n586), .Q(
        images_bus[111]) );
  dfcrq1 \images_bus_reg[326]  ( .D(n12927), .CP(clk), .CDN(n554), .Q(
        images_bus[326]) );
  dfcrq1 \images_bus_reg[402]  ( .D(n12851), .CP(clk), .CDN(n571), .Q(
        images_bus[402]) );
  dfcrq1 \images_bus_reg[14]  ( .D(n13239), .CP(clk), .CDN(n555), .Q(
        images_bus[14]) );
  dfcrq1 \images_bus_reg[291]  ( .D(n12962), .CP(clk), .CDN(n596), .Q(
        images_bus[291]) );
  dfcrq1 \images_bus_reg[157]  ( .D(n13096), .CP(clk), .CDN(n582), .Q(
        images_bus[157]) );
  dfcrq1 \images_bus_reg[64]  ( .D(n13189), .CP(clk), .CDN(n562), .Q(
        images_bus[64]) );
  dfcrq1 \images_bus_reg[257]  ( .D(n12996), .CP(clk), .CDN(n590), .Q(
        images_bus[257]) );
  dfcrq1 \images_bus_reg[139]  ( .D(n13114), .CP(clk), .CDN(n597), .Q(
        images_bus[139]) );
  dfcrq1 \images_bus_reg[62]  ( .D(n13191), .CP(clk), .CDN(n558), .Q(
        images_bus[62]) );
  dfcrq1 \images_bus_reg[223]  ( .D(n13030), .CP(clk), .CDN(n559), .Q(
        images_bus[223]) );
  dfcrq1 \images_bus_reg[146]  ( .D(n13107), .CP(clk), .CDN(n570), .Q(
        images_bus[146]) );
  dfcrq1 \images_bus_reg[76]  ( .D(n13177), .CP(clk), .CDN(n550), .Q(
        images_bus[76]) );
  dfcrq1 \images_bus_reg[239]  ( .D(n13014), .CP(clk), .CDN(n587), .Q(
        images_bus[239]) );
  dfcrq1 \images_bus_reg[46]  ( .D(n13207), .CP(clk), .CDN(n555), .Q(
        images_bus[46]) );
  dfcrq1 \images_bus_reg[105]  ( .D(n13148), .CP(clk), .CDN(n591), .Q(
        images_bus[105]) );
  dfcrq1 \images_bus_reg[404]  ( .D(n12849), .CP(clk), .CDN(n552), .Q(
        images_bus[404]) );
  dfcrq1 \images_bus_reg[11]  ( .D(n13242), .CP(clk), .CDN(n597), .Q(
        images_bus[11]) );
  dfcrq1 \images_bus_reg[184]  ( .D(n13069), .CP(clk), .CDN(n567), .Q(
        images_bus[184]) );
  dfcrq1 \images_bus_reg[51]  ( .D(n13202), .CP(clk), .CDN(n574), .Q(
        images_bus[51]) );
  dfcrq1 \images_bus_reg[32]  ( .D(n13221), .CP(clk), .CDN(n568), .Q(
        images_bus[32]) );
  dfcrq1 \images_bus_reg[85]  ( .D(n13168), .CP(clk), .CDN(n580), .Q(
        images_bus[85]) );
  dfcrq1 \images_bus_reg[117]  ( .D(n13136), .CP(clk), .CDN(n580), .Q(
        images_bus[117]) );
  dfcrq1 \images_bus_reg[70]  ( .D(n13183), .CP(clk), .CDN(n553), .Q(
        images_bus[70]) );
  dfcrq1 \images_bus_reg[182]  ( .D(n13071), .CP(clk), .CDN(n557), .Q(
        images_bus[182]) );
  dfcrq1 \images_bus_reg[120]  ( .D(n13133), .CP(clk), .CDN(n566), .Q(
        images_bus[120]) );
  dfcrq1 \images_bus_reg[300]  ( .D(n12953), .CP(clk), .CDN(n695), .Q(
        images_bus[300]) );
  dfcrq1 \images_bus_reg[332]  ( .D(n12921), .CP(clk), .CDN(n707), .Q(
        images_bus[332]) );
  dfcrq1 \images_bus_reg[66]  ( .D(n13187), .CP(clk), .CDN(n568), .Q(
        images_bus[66]) );
  dfcrq1 \images_bus_reg[358]  ( .D(n12895), .CP(clk), .CDN(n554), .Q(
        images_bus[358]) );
  dfcrq1 \images_bus_reg[71]  ( .D(n13182), .CP(clk), .CDN(n560), .Q(
        images_bus[71]) );
  dfcrq1 \images_bus_reg[40]  ( .D(n13213), .CP(clk), .CDN(n563), .Q(
        images_bus[40]) );
  dfcrq1 \images_bus_reg[123]  ( .D(n13130), .CP(clk), .CDN(n576), .Q(
        images_bus[123]) );
  dfcrq1 \images_bus_reg[438]  ( .D(n12815), .CP(clk), .CDN(n557), .Q(
        images_bus[438]) );
  dfcrq1 \images_bus_reg[322]  ( .D(n12931), .CP(clk), .CDN(n568), .Q(
        images_bus[322]) );
  dfcrq1 \images_bus_reg[371]  ( .D(n12882), .CP(clk), .CDN(n575), .Q(
        images_bus[371]) );
  dfcrq1 \images_bus_reg[368]  ( .D(n12885), .CP(clk), .CDN(n566), .Q(
        images_bus[368]) );
  dfcrq1 \images_bus_reg[374]  ( .D(n12879), .CP(clk), .CDN(n557), .Q(
        images_bus[374]) );
  dfcrq1 \images_bus_reg[89]  ( .D(n13164), .CP(clk), .CDN(n594), .Q(
        images_bus[89]) );
  dfcrq1 \images_bus_reg[262]  ( .D(n12991), .CP(clk), .CDN(n554), .Q(
        images_bus[262]) );
  dfcrq1 \images_bus_reg[415]  ( .D(n12838), .CP(clk), .CDN(n560), .Q(
        images_bus[415]) );
  dfcrq1 \images_bus_reg[310]  ( .D(n12943), .CP(clk), .CDN(n557), .Q(
        images_bus[310]) );
  dfcrq1 \images_bus_reg[297]  ( .D(n12956), .CP(clk), .CDN(n591), .Q(
        images_bus[297]) );
  dfcrq1 \images_bus_reg[334]  ( .D(n12919), .CP(clk), .CDN(n555), .Q(
        images_bus[334]) );
  dfcrq1 \images_bus_reg[69]  ( .D(n13184), .CP(clk), .CDN(n577), .Q(
        images_bus[69]) );
  dfcrq1 \images_bus_reg[47]  ( .D(n13206), .CP(clk), .CDN(n586), .Q(
        images_bus[47]) );
  dfcrq1 \images_bus_reg[340]  ( .D(n12913), .CP(clk), .CDN(n552), .Q(
        images_bus[340]) );
  dfcrq1 \images_bus_reg[299]  ( .D(n12954), .CP(clk), .CDN(n598), .Q(
        images_bus[299]) );
  dfcrq1 \images_bus_reg[345]  ( .D(n12908), .CP(clk), .CDN(n595), .Q(
        images_bus[345]) );
  dfcrq1 \images_bus_reg[439]  ( .D(n12814), .CP(clk), .CDN(n589), .Q(
        images_bus[439]) );
  dfcrq1 \images_bus_reg[360]  ( .D(n12893), .CP(clk), .CDN(n564), .Q(
        images_bus[360]) );
  dfcrq1 \images_bus_reg[362]  ( .D(n12891), .CP(clk), .CDN(n570), .Q(
        images_bus[362]) );
  dfcrq1 \images_bus_reg[373]  ( .D(n12880), .CP(clk), .CDN(n581), .Q(
        images_bus[373]) );
  dfcrq1 \images_bus_reg[136]  ( .D(n13117), .CP(clk), .CDN(n563), .Q(
        images_bus[136]) );
  dfcrq1 \images_bus_reg[86]  ( .D(n13167), .CP(clk), .CDN(n556), .Q(
        images_bus[86]) );
  dfcrq1 \images_bus_reg[273]  ( .D(n12980), .CP(clk), .CDN(n593), .Q(
        images_bus[273]) );
  dfcrq1 \images_bus_reg[305]  ( .D(n12948), .CP(clk), .CDN(n593), .Q(
        images_bus[305]) );
  dfcrq1 \images_bus_reg[20]  ( .D(n13233), .CP(clk), .CDN(n551), .Q(
        images_bus[20]) );
  dfcrq1 \images_bus_reg[207]  ( .D(n13046), .CP(clk), .CDN(n586), .Q(
        images_bus[207]) );
  dfcrq1 \images_bus_reg[348]  ( .D(n12905), .CP(clk), .CDN(n553), .Q(
        images_bus[348]) );
  dfcrq1 \images_bus_reg[359]  ( .D(n12894), .CP(clk), .CDN(n561), .Q(
        images_bus[359]) );
  dfcrq1 \images_bus_reg[400]  ( .D(n12853), .CP(clk), .CDN(n566), .Q(
        images_bus[400]) );
  dfcrq1 \images_bus_reg[222]  ( .D(n13031), .CP(clk), .CDN(n558), .Q(
        images_bus[222]) );
  dfcrq1 \images_bus_reg[168]  ( .D(n13085), .CP(clk), .CDN(n564), .Q(
        images_bus[168]) );
  dfcrq1 \images_bus_reg[302]  ( .D(n12951), .CP(clk), .CDN(n555), .Q(
        images_bus[302]) );
  dfcrq1 \images_bus_reg[366]  ( .D(n12887), .CP(clk), .CDN(n556), .Q(
        images_bus[366]) );
  dfcrq1 \images_bus_reg[270]  ( .D(n12983), .CP(clk), .CDN(n555), .Q(
        images_bus[270]) );
  dfcrq1 \images_bus_reg[60]  ( .D(n13193), .CP(clk), .CDN(n552), .Q(
        images_bus[60]) );
  dfcrq1 \images_bus_reg[77]  ( .D(n13176), .CP(clk), .CDN(n579), .Q(
        images_bus[77]) );
  dfcrq1 \images_bus_reg[103]  ( .D(n13150), .CP(clk), .CDN(n560), .Q(
        images_bus[103]) );
  dfcrq1 \images_bus_reg[121]  ( .D(n13132), .CP(clk), .CDN(n594), .Q(
        images_bus[121]) );
  dfcrq1 \images_bus_reg[125]  ( .D(n13128), .CP(clk), .CDN(n582), .Q(
        images_bus[125]) );
  dfcrq1 \images_bus_reg[331]  ( .D(n12922), .CP(clk), .CDN(n598), .Q(
        images_bus[331]) );
  dfcrq1 \images_bus_reg[288]  ( .D(n12965), .CP(clk), .CDN(n562), .Q(
        images_bus[288]) );
  dfcrq1 \images_bus_reg[41]  ( .D(n13212), .CP(clk), .CDN(n591), .Q(
        images_bus[41]) );
  dfcrq1 \images_bus_reg[17]  ( .D(n13236), .CP(clk), .CDN(n592), .Q(
        images_bus[17]) );
  dfcrq1 \images_bus_reg[399]  ( .D(n12854), .CP(clk), .CDN(n587), .Q(
        images_bus[399]) );
  dfcrq1 \images_bus_reg[479]  ( .D(n12774), .CP(clk), .CDN(n560), .Q(
        images_bus[479]) );
  dfcrq1 \images_bus_reg[28]  ( .D(n13225), .CP(clk), .CDN(n552), .Q(
        images_bus[28]) );
  dfcrq1 \images_bus_reg[293]  ( .D(n12960), .CP(clk), .CDN(n578), .Q(
        images_bus[293]) );
  dfcrq1 \images_bus_reg[93]  ( .D(n13160), .CP(clk), .CDN(n582), .Q(
        images_bus[93]) );
  dfcrq1 \images_bus_reg[12]  ( .D(n13241), .CP(clk), .CDN(n574), .Q(
        images_bus[12]) );
  dfcrq1 \images_bus_reg[364]  ( .D(n12889), .CP(clk), .CDN(n551), .Q(
        images_bus[364]) );
  dfcrq1 \images_bus_reg[25]  ( .D(n13228), .CP(clk), .CDN(n594), .Q(
        images_bus[25]) );
  dfcrq1 \images_bus_reg[48]  ( .D(n13205), .CP(clk), .CDN(n565), .Q(
        images_bus[48]) );
  dfcrq1 \images_bus_reg[106]  ( .D(n13147), .CP(clk), .CDN(n569), .Q(
        images_bus[106]) );
  dfcrq1 \images_bus_reg[333]  ( .D(n12920), .CP(clk), .CDN(n580), .Q(
        images_bus[333]) );
  dfcrq1 \images_bus_reg[407]  ( .D(n12846), .CP(clk), .CDN(n589), .Q(
        images_bus[407]) );
  dfcrq1 \images_bus_reg[152]  ( .D(n13101), .CP(clk), .CDN(n566), .Q(
        images_bus[152]) );
  dfcrq1 \images_bus_reg[339]  ( .D(n12914), .CP(clk), .CDN(n575), .Q(
        images_bus[339]) );
  dfcrq1 \images_bus_reg[328]  ( .D(n12925), .CP(clk), .CDN(n564), .Q(
        images_bus[328]) );
  dfcrq1 \images_bus_reg[256]  ( .D(n12997), .CP(clk), .CDN(n562), .Q(
        images_bus[256]) );
  dfcrq1 \images_bus_reg[44]  ( .D(n13209), .CP(clk), .CDN(n556), .Q(
        images_bus[44]) );
  dfcrq1 \images_bus_reg[265]  ( .D(n12988), .CP(clk), .CDN(n591), .Q(
        images_bus[265]) );
  dfcrq1 \images_bus_reg[79]  ( .D(n13174), .CP(clk), .CDN(n586), .Q(
        images_bus[79]) );
  dfcrq1 \images_bus_reg[87]  ( .D(n13166), .CP(clk), .CDN(n588), .Q(
        images_bus[87]) );
  dfcrq1 \images_bus_reg[159]  ( .D(n13094), .CP(clk), .CDN(n559), .Q(
        images_bus[159]) );
  dfcrq1 \images_bus_reg[54]  ( .D(n13199), .CP(clk), .CDN(n556), .Q(
        images_bus[54]) );
  dfcrq1 \images_bus_reg[376]  ( .D(n12877), .CP(clk), .CDN(n567), .Q(
        images_bus[376]) );
  dfcrq1 \images_bus_reg[6]  ( .D(n13247), .CP(clk), .CDN(n553), .Q(
        images_bus[6]) );
  dfcrq1 \images_bus_reg[363]  ( .D(n12890), .CP(clk), .CDN(n580), .Q(
        images_bus[363]) );
  dfcrq1 \images_bus_reg[323]  ( .D(n12930), .CP(clk), .CDN(n596), .Q(
        images_bus[323]) );
  dfcrq1 \images_bus_reg[306]  ( .D(n12947), .CP(clk), .CDN(n571), .Q(
        images_bus[306]) );
  dfcrq1 \images_bus_reg[13]  ( .D(n13240), .CP(clk), .CDN(n579), .Q(
        images_bus[13]) );
  dfcrq1 \images_bus_reg[263]  ( .D(n12990), .CP(clk), .CDN(n561), .Q(
        images_bus[263]) );
  dfcrq1 \images_bus_reg[154]  ( .D(n13099), .CP(clk), .CDN(n572), .Q(
        images_bus[154]) );
  dfcrq1 \images_bus_reg[383]  ( .D(n12870), .CP(clk), .CDN(n560), .Q(
        images_bus[383]) );
  dfcrq1 \images_bus_reg[95]  ( .D(n13158), .CP(clk), .CDN(n559), .Q(
        images_bus[95]) );
  dfcrq1 \images_bus_reg[143]  ( .D(n13110), .CP(clk), .CDN(n586), .Q(
        images_bus[143]) );
  dfcrq1 \images_bus_reg[122]  ( .D(n13131), .CP(clk), .CDN(n571), .Q(
        images_bus[122]) );
  dfcrq1 \images_bus_reg[301]  ( .D(n12952), .CP(clk), .CDN(n580), .Q(
        images_bus[301]) );
  dfcrq1 \images_bus_reg[8]  ( .D(n13245), .CP(clk), .CDN(n563), .Q(
        images_bus[8]) );
  dfcrq1 \images_bus_reg[382]  ( .D(n12871), .CP(clk), .CDN(n558), .Q(
        images_bus[382]) );
  dfcrq1 \images_bus_reg[59]  ( .D(n13194), .CP(clk), .CDN(n576), .Q(
        images_bus[59]) );
  dfcrq1 \images_bus_reg[29]  ( .D(n13224), .CP(clk), .CDN(n582), .Q(
        images_bus[29]) );
  dfcrq1 \images_bus_reg[126]  ( .D(n13127), .CP(clk), .CDN(n558), .Q(
        images_bus[126]) );
  dfcrq1 \images_bus_reg[336]  ( .D(n12917), .CP(clk), .CDN(n566), .Q(
        images_bus[336]) );
  dfcrq1 \images_bus_reg[7]  ( .D(n13246), .CP(clk), .CDN(n560), .Q(
        images_bus[7]) );
  dfcrq1 \images_bus_reg[258]  ( .D(n12995), .CP(clk), .CDN(n568), .Q(
        images_bus[258]) );
  dfcrq1 \images_bus_reg[330]  ( .D(n12923), .CP(clk), .CDN(n569), .Q(
        images_bus[330]) );
  dfcrq1 \images_bus_reg[381]  ( .D(n12872), .CP(clk), .CDN(n583), .Q(
        images_bus[381]) );
  dfcrq1 \images_bus_reg[61]  ( .D(n13192), .CP(clk), .CDN(n582), .Q(
        images_bus[61]) );
  dfcrq1 \images_bus_reg[367]  ( .D(n12886), .CP(clk), .CDN(n587), .Q(
        images_bus[367]) );
  dfcrq1 \images_bus_reg[175]  ( .D(n13078), .CP(clk), .CDN(n586), .Q(
        images_bus[175]) );
  dfcrq1 \images_bus_reg[278]  ( .D(n12975), .CP(clk), .CDN(n557), .Q(
        images_bus[278]) );
  dfcrq1 \images_bus_reg[335]  ( .D(n12918), .CP(clk), .CDN(n587), .Q(
        images_bus[335]) );
  dfcrq1 \images_bus_reg[296]  ( .D(n12957), .CP(clk), .CDN(n564), .Q(
        images_bus[296]) );
  dfcrq1 \images_bus_reg[349]  ( .D(n12904), .CP(clk), .CDN(n583), .Q(
        images_bus[349]) );
  dfcrq1 \images_bus_reg[21]  ( .D(n13232), .CP(clk), .CDN(n580), .Q(
        images_bus[21]) );
  dfcrq1 \images_bus_reg[74]  ( .D(n13179), .CP(clk), .CDN(n569), .Q(
        images_bus[74]) );
  dfcrq1 \images_bus_reg[343]  ( .D(n12910), .CP(clk), .CDN(n588), .Q(
        images_bus[343]) );
  dfcrq1 \images_bus_reg[88]  ( .D(n13165), .CP(clk), .CDN(n566), .Q(
        images_bus[88]) );
  dfcrq1 \images_bus_reg[23]  ( .D(n13230), .CP(clk), .CDN(n587), .Q(
        images_bus[23]) );
  dfcrq1 \images_bus_reg[82]  ( .D(n13171), .CP(clk), .CDN(n570), .Q(
        images_bus[82]) );
  dfcrq1 \images_bus_reg[380]  ( .D(n12873), .CP(clk), .CDN(n553), .Q(
        images_bus[380]) );
  dfcrq1 \images_bus_reg[45]  ( .D(n13208), .CP(clk), .CDN(n579), .Q(
        images_bus[45]) );
  dfcrq1 \images_bus_reg[277]  ( .D(n12976), .CP(clk), .CDN(n581), .Q(
        images_bus[277]) );
  dfcrq1 \images_bus_reg[324]  ( .D(n12929), .CP(clk), .CDN(n573), .Q(
        images_bus[324]) );
  dfcrq1 \images_bus_reg[269]  ( .D(n12984), .CP(clk), .CDN(n579), .Q(
        images_bus[269]) );
  dfcrq1 \images_bus_reg[281]  ( .D(n12972), .CP(clk), .CDN(n594), .Q(
        images_bus[281]) );
  dfcrq1 \images_bus_reg[42]  ( .D(n13211), .CP(clk), .CDN(n569), .Q(
        images_bus[42]) );
  dfcrq1 \images_bus_reg[309]  ( .D(n12944), .CP(clk), .CDN(n581), .Q(
        images_bus[309]) );
  dfcrq1 \compare_image_index_reg[7]  ( .D(n12196), .CP(clk), .CDN(n585), .Q(
        N3181) );
  dfcrq1 \images_bus_reg[304]  ( .D(n12949), .CP(clk), .CDN(n565), .Q(
        images_bus[304]) );
  dfcrq1 \images_bus_reg[56]  ( .D(n13197), .CP(clk), .CDN(n566), .Q(
        images_bus[56]) );
  dfcrq1 \images_bus_reg[316]  ( .D(n12937), .CP(clk), .CDN(n553), .Q(
        images_bus[316]) );
  dfcrq1 \images_bus_reg[94]  ( .D(n13159), .CP(clk), .CDN(n558), .Q(
        images_bus[94]) );
  dfcrq1 \images_bus_reg[57]  ( .D(n13196), .CP(clk), .CDN(n594), .Q(
        images_bus[57]) );
  dfcrq1 \images_bus_reg[341]  ( .D(n12912), .CP(clk), .CDN(n581), .Q(
        images_bus[341]) );
  dfcrq1 \images_bus_reg[259]  ( .D(n12994), .CP(clk), .CDN(n596), .Q(
        images_bus[259]) );
  dfcrq1 \images_bus_reg[30]  ( .D(n13223), .CP(clk), .CDN(n557), .Q(
        images_bus[30]) );
  dfcrq1 \images_bus_reg[22]  ( .D(n13231), .CP(clk), .CDN(n556), .Q(
        images_bus[22]) );
  dfcrq1 \images_bus_reg[276]  ( .D(n12977), .CP(clk), .CDN(n551), .Q(
        images_bus[276]) );
  dfcrq1 \images_bus_reg[91]  ( .D(n13162), .CP(clk), .CDN(n576), .Q(
        images_bus[91]) );
  dfcrq1 \images_bus_reg[351]  ( .D(n12902), .CP(clk), .CDN(n560), .Q(
        images_bus[351]) );
  dfcrq1 \images_bus_reg[16]  ( .D(n13237), .CP(clk), .CDN(n565), .Q(
        images_bus[16]) );
  dfcrq1 \images_bus_reg[279]  ( .D(n12974), .CP(clk), .CDN(n588), .Q(
        images_bus[279]) );
  dfcrq1 \images_bus_reg[275]  ( .D(n12978), .CP(clk), .CDN(n575), .Q(
        images_bus[275]) );
  dfcrq1 \images_bus_reg[298]  ( .D(n12955), .CP(clk), .CDN(n569), .Q(
        images_bus[298]) );
  dfcrq1 \images_bus_reg[313]  ( .D(n12940), .CP(clk), .CDN(n595), .Q(
        images_bus[313]) );
  dfcrq1 \images_bus_reg[327]  ( .D(n12926), .CP(clk), .CDN(n561), .Q(
        images_bus[327]) );
  dfcrq1 \images_bus_reg[272]  ( .D(n12981), .CP(clk), .CDN(n565), .Q(
        images_bus[272]) );
  dfcrq1 \images_bus_reg[344]  ( .D(n12909), .CP(clk), .CDN(n567), .Q(
        images_bus[344]) );
  dfcrq1 \images_bus_reg[379]  ( .D(n12874), .CP(clk), .CDN(n577), .Q(
        images_bus[379]) );
  dfcrq1 \images_bus_reg[338]  ( .D(n12915), .CP(clk), .CDN(n571), .Q(
        images_bus[338]) );
  dfcrq1 \images_bus_reg[318]  ( .D(n12935), .CP(clk), .CDN(n558), .Q(
        images_bus[318]) );
  dfcrq1 \images_bus_reg[63]  ( .D(n13190), .CP(clk), .CDN(n559), .Q(
        images_bus[63]) );
  dfcrq1 \images_bus_reg[19]  ( .D(n13234), .CP(clk), .CDN(n574), .Q(
        images_bus[19]) );
  dfcrq1 \images_bus_reg[24]  ( .D(n13229), .CP(clk), .CDN(n566), .Q(
        images_bus[24]) );
  dfcrq1 \images_bus_reg[15]  ( .D(n13238), .CP(clk), .CDN(n586), .Q(
        images_bus[15]) );
  dfcrq1 \images_bus_reg[31]  ( .D(n13222), .CP(clk), .CDN(n559), .Q(
        images_bus[31]) );
  dfcrq1 \images_bus_reg[295]  ( .D(n12958), .CP(clk), .CDN(n561), .Q(
        images_bus[295]) );
  dfcrq1 \images_bus_reg[267]  ( .D(n12986), .CP(clk), .CDN(n598), .Q(
        images_bus[267]) );
  dfcrq1 \images_bus_reg[312]  ( .D(n12941), .CP(clk), .CDN(n567), .Q(
        images_bus[312]) );
  dfcrq1 \images_bus_reg[268]  ( .D(n12985), .CP(clk), .CDN(n550), .Q(
        images_bus[268]) );
  dfcrq1 \images_bus_reg[350]  ( .D(n12903), .CP(clk), .CDN(n558), .Q(
        images_bus[350]) );
  dfcrq1 \images_bus_reg[18]  ( .D(n13235), .CP(clk), .CDN(n570), .Q(
        images_bus[18]) );
  dfcrq1 \images_bus_reg[58]  ( .D(n13195), .CP(clk), .CDN(n571), .Q(
        images_bus[58]) );
  dfcrq1 \images_bus_reg[26]  ( .D(n13227), .CP(clk), .CDN(n571), .Q(
        images_bus[26]) );
  dfcrq1 \images_bus_reg[127]  ( .D(n13126), .CP(clk), .CDN(n559), .Q(
        images_bus[127]) );
  dfcrq1 \images_bus_reg[375]  ( .D(n12878), .CP(clk), .CDN(n589), .Q(
        images_bus[375]) );
  dfcrq1 \images_bus_reg[271]  ( .D(n12982), .CP(clk), .CDN(n587), .Q(
        images_bus[271]) );
  dfcrq1 \images_bus_reg[119]  ( .D(n13134), .CP(clk), .CDN(n588), .Q(
        images_bus[119]) );
  dfcrq1 \images_bus_reg[104]  ( .D(n13149), .CP(clk), .CDN(n563), .Q(
        images_bus[104]) );
  dfcrq1 \images_bus_reg[347]  ( .D(n12906), .CP(clk), .CDN(n577), .Q(
        images_bus[347]) );
  dfcrq1 \images_bus_reg[285]  ( .D(n12968), .CP(clk), .CDN(n582), .Q(
        images_bus[285]) );
  dfcrq1 \images_bus_reg[314]  ( .D(n12939), .CP(clk), .CDN(n572), .Q(
        images_bus[314]) );
  dfcrq1 \images_bus_reg[55]  ( .D(n13198), .CP(clk), .CDN(n588), .Q(
        images_bus[55]) );
  dfcrq1 \images_bus_reg[266]  ( .D(n12987), .CP(clk), .CDN(n569), .Q(
        images_bus[266]) );
  dfcrq1 \images_bus_reg[307]  ( .D(n12946), .CP(clk), .CDN(n575), .Q(
        images_bus[307]) );
  dfcrq1 \images_bus_reg[27]  ( .D(n13226), .CP(clk), .CDN(n576), .Q(
        images_bus[27]) );
  dfcrq1 \images_bus_reg[286]  ( .D(n12967), .CP(clk), .CDN(n558), .Q(
        images_bus[286]) );
  dfcrq1 \images_bus_reg[315]  ( .D(n12938), .CP(clk), .CDN(n576), .Q(
        images_bus[315]) );
  dfcrq1 \images_bus_reg[280]  ( .D(n12973), .CP(clk), .CDN(n567), .Q(
        images_bus[280]) );
  dfcrq1 \images_bus_reg[282]  ( .D(n12971), .CP(clk), .CDN(n572), .Q(
        images_bus[282]) );
  dfcrq1 \images_bus_reg[287]  ( .D(n12966), .CP(clk), .CDN(n559), .Q(
        images_bus[287]) );
  dfcrq1 \images_bus_reg[311]  ( .D(n12942), .CP(clk), .CDN(n588), .Q(
        images_bus[311]) );
  dfcrq1 \images_bus_reg[2]  ( .D(n13251), .CP(clk), .CDN(n568), .Q(
        images_bus[2]) );
  dfcrq1 \images_bus_reg[317]  ( .D(n12936), .CP(clk), .CDN(n583), .Q(
        images_bus[317]) );
  dfcrq1 \images_bus_reg[274]  ( .D(n12979), .CP(clk), .CDN(n571), .Q(
        images_bus[274]) );
  dfcrq1 \images_bus_reg[319]  ( .D(n12934), .CP(clk), .CDN(n560), .Q(
        images_bus[319]) );
  dfcrq1 \images_bus_reg[264]  ( .D(n12989), .CP(clk), .CDN(n564), .Q(
        images_bus[264]) );
  dfcrq1 \images_bus_reg[346]  ( .D(n12907), .CP(clk), .CDN(n572), .Q(
        images_bus[346]) );
  dfcrq1 \images_bus_reg[303]  ( .D(n12950), .CP(clk), .CDN(n587), .Q(
        images_bus[303]) );
  dfcrq1 \count_image_reg[3]  ( .D(n12738), .CP(clk), .CDN(n584), .Q(
        count_image[3]) );
  dfcrq1 \count_image_reg[7]  ( .D(n12734), .CP(clk), .CDN(n584), .Q(
        count_image[7]) );
  dfcrq1 \compare_image_index_reg[3]  ( .D(n12192), .CP(clk), .CDN(n585), .Q(
        N3975) );
  dfcrq1 \compare_image_index_reg[5]  ( .D(n12194), .CP(clk), .CDN(n585), .Q(
        N3179) );
  dfcrq1 \compare_image_index_reg[4]  ( .D(n12193), .CP(clk), .CDN(n585), .Q(
        N3976) );
  dfcrq1 \compare_image_index_reg[0]  ( .D(n12201), .CP(clk), .CDN(n574), .Q(
        N3972) );
  dfcrq1 \compare_image_index_reg[1]  ( .D(n12190), .CP(clk), .CDN(n585), .Q(
        N3973) );
  dfcrq1 \compare_image_index_reg[2]  ( .D(n12191), .CP(clk), .CDN(n585), .Q(
        N3974) );
  dfnrq1 \reorder_A2_reg[8]  ( .D(n12101), .CP(clk), .Q(reorder_A2[8]) );
  dfnrq1 \reorder_A2_reg[0]  ( .D(n12093), .CP(clk), .Q(reorder_A2[0]) );
  dfnrq1 \reorder_A2_reg[2]  ( .D(n12095), .CP(clk), .Q(reorder_A2[2]) );
  dfnrq1 \reorder_A2_reg[1]  ( .D(n12094), .CP(clk), .Q(reorder_A2[1]) );
  dfnrq1 \reorder_A2_reg[11]  ( .D(n12104), .CP(clk), .Q(reorder_A2[11]) );
  dfnrq1 \reorder_A2_reg[10]  ( .D(n12103), .CP(clk), .Q(reorder_A2[10]) );
  dfnrq1 \reorder_A2_reg[9]  ( .D(n12102), .CP(clk), .Q(reorder_A2[9]) );
  dfnrq1 \reorder_A2_reg[7]  ( .D(n12100), .CP(clk), .Q(reorder_A2[7]) );
  dfnrq1 \reorder_A2_reg[6]  ( .D(n12099), .CP(clk), .Q(reorder_A2[6]) );
  dfnrq1 \reorder_A2_reg[5]  ( .D(n12098), .CP(clk), .Q(reorder_A2[5]) );
  dfnrq1 \reorder_A2_reg[4]  ( .D(n12097), .CP(clk), .Q(reorder_A2[4]) );
  dfnrq1 \reorder_A2_reg[3]  ( .D(n12096), .CP(clk), .Q(reorder_A2[3]) );
  dfnrq1 \reorder_A1_reg[2]  ( .D(n12107), .CP(clk), .Q(reorder_A1[2]) );
  dfnrq1 \reorder_A1_reg[1]  ( .D(n12106), .CP(clk), .Q(reorder_A1[1]) );
  dfnrq1 \reorder_A1_reg[0]  ( .D(n12105), .CP(clk), .Q(reorder_A1[0]) );
  dfnrq1 \reorder_A1_reg[11]  ( .D(n12116), .CP(clk), .Q(reorder_A1[11]) );
  dfnrq1 \reorder_A1_reg[10]  ( .D(n12115), .CP(clk), .Q(reorder_A1[10]) );
  dfnrq1 \reorder_A1_reg[9]  ( .D(n12114), .CP(clk), .Q(reorder_A1[9]) );
  dfnrq1 \reorder_A1_reg[8]  ( .D(n12113), .CP(clk), .Q(reorder_A1[8]) );
  dfnrq1 \reorder_A1_reg[7]  ( .D(n12112), .CP(clk), .Q(reorder_A1[7]) );
  dfnrq1 \reorder_A1_reg[6]  ( .D(n12111), .CP(clk), .Q(reorder_A1[6]) );
  dfnrq1 \reorder_A1_reg[5]  ( .D(n12110), .CP(clk), .Q(reorder_A1[5]) );
  dfnrq1 \reorder_A1_reg[4]  ( .D(n12109), .CP(clk), .Q(reorder_A1[4]) );
  dfnrq1 \reorder_A1_reg[3]  ( .D(n12108), .CP(clk), .Q(reorder_A1[3]) );
  aoim21d1 U2307 ( .B1(n4337), .B2(1'b0), .A(n2768), .ZN(n4363) );
  aoim21d1 U2272 ( .B1(1'b0), .B2(n4329), .A(n2768), .ZN(n4360) );
  aoim21d1 U2377 ( .B1(n4345), .B2(1'b0), .A(n2768), .ZN(n4370) );
  aoim21d1 U2342 ( .B1(1'b0), .B2(n4337), .A(n2768), .ZN(n4367) );
  aoim21d1 U2474 ( .B1(1'b0), .B2(n4345), .A(n2768), .ZN(n4372) );
  aoim21d1 U2483 ( .B1(n2781), .B2(1'b0), .A(n2768), .ZN(n4356) );
  aoim21d1 U2239 ( .B1(1'b0), .B2(n4329), .A(n2768), .ZN(n4359) );
  aoim21d1 U2173 ( .B1(n2781), .B2(1'b0), .A(n2768), .ZN(n4353) );
  ad01d0 \add_0_root_add_1_root_add_130_3/U1_4  ( .A(N3973), .B(1'b0), .CI(
        \add_0_root_add_1_root_add_130_3/carry[4] ), .CO(
        \add_0_root_add_1_root_add_130_3/carry[5] ), .S(N4689) );
  ad01d0 \add_0_root_add_1_root_add_98_3/U1_4  ( .A(
        \add_0_root_add_1_root_add_98_3/A[4] ), .B(1'b0), .CI(
        \add_0_root_add_1_root_add_98_3/carry[4] ), .CO(
        \add_0_root_add_1_root_add_98_3/carry[5] ), .S(N3880) );
  nr04d1 U2344 ( .A1(n2789), .A2(1'b0), .A3(N3877), .A4(N3855), .ZN(n4337) );
  oai222d1 U2306 ( .A1(n7558), .A2(1'b1), .B1(n12628), .B2(n756), .C1(n7408), 
        .C2(n750), .ZN(n13695) );
  oai222d1 U2305 ( .A1(n7514), .A2(1'b1), .B1(n12627), .B2(n756), .C1(n7377), 
        .C2(n750), .ZN(n13694) );
  oai222d1 U2304 ( .A1(n7448), .A2(1'b1), .B1(n12626), .B2(n756), .C1(n7318), 
        .C2(n750), .ZN(n13693) );
  oai222d1 U2303 ( .A1(n7438), .A2(1'b1), .B1(n12625), .B2(n756), .C1(n7297), 
        .C2(n750), .ZN(n13692) );
  oai222d1 U2302 ( .A1(n7432), .A2(1'b1), .B1(n12624), .B2(n756), .C1(n7293), 
        .C2(n750), .ZN(n13691) );
  oai222d1 U2301 ( .A1(n7425), .A2(1'b1), .B1(n12623), .B2(n756), .C1(n7288), 
        .C2(n749), .ZN(n13690) );
  oai222d1 U2300 ( .A1(n7424), .A2(1'b1), .B1(n12622), .B2(n756), .C1(n7278), 
        .C2(n749), .ZN(n13689) );
  oai222d1 U2299 ( .A1(n7415), .A2(1'b1), .B1(n12621), .B2(n756), .C1(n7271), 
        .C2(n749), .ZN(n13688) );
  oai222d1 U2298 ( .A1(n7414), .A2(1'b1), .B1(n12620), .B2(n756), .C1(n7265), 
        .C2(n749), .ZN(n13687) );
  oai222d1 U2297 ( .A1(n7412), .A2(1'b1), .B1(n12619), .B2(n757), .C1(n7261), 
        .C2(n749), .ZN(n13686) );
  oai222d1 U2296 ( .A1(n7553), .A2(1'b1), .B1(n12618), .B2(n757), .C1(n7405), 
        .C2(n749), .ZN(n13685) );
  oai222d1 U2295 ( .A1(n7552), .A2(1'b1), .B1(n12617), .B2(n757), .C1(n7403), 
        .C2(n749), .ZN(n13684) );
  oai222d1 U2294 ( .A1(n7549), .A2(1'b1), .B1(n12616), .B2(n757), .C1(n7402), 
        .C2(n749), .ZN(n13683) );
  oai222d1 U2293 ( .A1(n7542), .A2(1'b1), .B1(n12615), .B2(n757), .C1(n7399), 
        .C2(n749), .ZN(n13682) );
  oai222d1 U2292 ( .A1(n7538), .A2(1'b1), .B1(n12614), .B2(n757), .C1(n7398), 
        .C2(n748), .ZN(n13681) );
  oai222d1 U2291 ( .A1(n7531), .A2(1'b1), .B1(n12613), .B2(n757), .C1(n7397), 
        .C2(n748), .ZN(n13680) );
  oai222d1 U2290 ( .A1(n7525), .A2(1'b1), .B1(n12612), .B2(n757), .C1(n7390), 
        .C2(n748), .ZN(n13679) );
  oai222d1 U2289 ( .A1(n7524), .A2(1'b1), .B1(n12611), .B2(n757), .C1(n7387), 
        .C2(n748), .ZN(n13678) );
  oai222d1 U2288 ( .A1(n7520), .A2(1'b1), .B1(n12610), .B2(n758), .C1(n7380), 
        .C2(n748), .ZN(n13677) );
  oai222d1 U2287 ( .A1(n7519), .A2(1'b1), .B1(n12609), .B2(n758), .C1(n7379), 
        .C2(n748), .ZN(n13676) );
  oai222d1 U2286 ( .A1(n7510), .A2(1'b1), .B1(n12608), .B2(n758), .C1(n7372), 
        .C2(n748), .ZN(n13675) );
  oai222d1 U2285 ( .A1(n7503), .A2(1'b1), .B1(n12607), .B2(n758), .C1(n7371), 
        .C2(n748), .ZN(n13674) );
  oai222d1 U2284 ( .A1(n7497), .A2(1'b1), .B1(n12606), .B2(n758), .C1(n7365), 
        .C2(n748), .ZN(n13673) );
  oai222d1 U2283 ( .A1(n7482), .A2(1'b1), .B1(n12605), .B2(n758), .C1(n7363), 
        .C2(n747), .ZN(n13672) );
  oai222d1 U2282 ( .A1(n7476), .A2(1'b1), .B1(n12604), .B2(n758), .C1(n7361), 
        .C2(n747), .ZN(n13671) );
  oai222d1 U2281 ( .A1(n7470), .A2(1'b1), .B1(n12603), .B2(n758), .C1(n7355), 
        .C2(n747), .ZN(n13670) );
  oai222d1 U2280 ( .A1(n7467), .A2(1'b1), .B1(n12602), .B2(n758), .C1(n7348), 
        .C2(n747), .ZN(n13669) );
  oai222d1 U2279 ( .A1(n7465), .A2(1'b1), .B1(n12601), .B2(n759), .C1(n7342), 
        .C2(n747), .ZN(n13668) );
  oai222d1 U2278 ( .A1(n7451), .A2(1'b1), .B1(n12600), .B2(n759), .C1(n7325), 
        .C2(n747), .ZN(n13667) );
  oai222d1 U2277 ( .A1(n7449), .A2(1'b1), .B1(n12599), .B2(n759), .C1(n7322), 
        .C2(n747), .ZN(n13666) );
  oai222d1 U2276 ( .A1(n7445), .A2(1'b1), .B1(n12598), .B2(n759), .C1(n7312), 
        .C2(n747), .ZN(n13665) );
  oai222d1 U2275 ( .A1(n7441), .A2(1'b1), .B1(n12597), .B2(n759), .C1(n7307), 
        .C2(n747), .ZN(n13664) );
  oai222d1 U2271 ( .A1(n7558), .A2(n782), .B1(n12596), .B2(n769), .C1(n7408), 
        .C2(1'b1), .ZN(n13663) );
  oai222d1 U2270 ( .A1(n7514), .A2(n782), .B1(n12595), .B2(n769), .C1(n7377), 
        .C2(1'b1), .ZN(n13662) );
  oai222d1 U2269 ( .A1(n7448), .A2(n782), .B1(n12594), .B2(n769), .C1(n7318), 
        .C2(1'b1), .ZN(n13661) );
  oai222d1 U2268 ( .A1(n7438), .A2(n782), .B1(n12593), .B2(n769), .C1(n7297), 
        .C2(1'b1), .ZN(n13660) );
  oai222d1 U2267 ( .A1(n7432), .A2(n782), .B1(n12592), .B2(n769), .C1(n7293), 
        .C2(1'b1), .ZN(n13659) );
  oai222d1 U2266 ( .A1(n7425), .A2(n782), .B1(n12591), .B2(n769), .C1(n7288), 
        .C2(1'b1), .ZN(n13658) );
  oai222d1 U2265 ( .A1(n7424), .A2(n782), .B1(n12590), .B2(n769), .C1(n7278), 
        .C2(1'b1), .ZN(n13657) );
  oai222d1 U2264 ( .A1(n7415), .A2(n782), .B1(n12589), .B2(n769), .C1(n7271), 
        .C2(1'b1), .ZN(n13656) );
  oai222d1 U2263 ( .A1(n7414), .A2(n782), .B1(n12588), .B2(n769), .C1(n7265), 
        .C2(1'b1), .ZN(n13655) );
  oai222d1 U2262 ( .A1(n7412), .A2(n783), .B1(n12587), .B2(n770), .C1(n7261), 
        .C2(1'b1), .ZN(n13654) );
  oai222d1 U2261 ( .A1(n7553), .A2(n783), .B1(n12586), .B2(n770), .C1(n7405), 
        .C2(1'b1), .ZN(n13653) );
  oai222d1 U2260 ( .A1(n7552), .A2(n783), .B1(n12585), .B2(n770), .C1(n7403), 
        .C2(1'b1), .ZN(n13652) );
  oai222d1 U2259 ( .A1(n7549), .A2(n783), .B1(n12584), .B2(n770), .C1(n7402), 
        .C2(1'b1), .ZN(n13651) );
  oai222d1 U2258 ( .A1(n7542), .A2(n783), .B1(n12583), .B2(n770), .C1(n7399), 
        .C2(1'b1), .ZN(n13650) );
  oai222d1 U2257 ( .A1(n7538), .A2(n783), .B1(n12582), .B2(n770), .C1(n7398), 
        .C2(1'b1), .ZN(n13649) );
  oai222d1 U2256 ( .A1(n7531), .A2(n783), .B1(n12581), .B2(n770), .C1(n7397), 
        .C2(1'b1), .ZN(n13648) );
  oai222d1 U2255 ( .A1(n7525), .A2(n783), .B1(n12580), .B2(n770), .C1(n7390), 
        .C2(1'b1), .ZN(n13647) );
  oai222d1 U2254 ( .A1(n7524), .A2(n783), .B1(n12579), .B2(n770), .C1(n7387), 
        .C2(1'b1), .ZN(n13646) );
  oai222d1 U2253 ( .A1(n7520), .A2(n784), .B1(n12578), .B2(n771), .C1(n7380), 
        .C2(1'b1), .ZN(n13645) );
  oai222d1 U2252 ( .A1(n7519), .A2(n784), .B1(n12577), .B2(n771), .C1(n7379), 
        .C2(1'b1), .ZN(n13644) );
  oai222d1 U2251 ( .A1(n7510), .A2(n784), .B1(n12576), .B2(n771), .C1(n7372), 
        .C2(1'b1), .ZN(n13643) );
  oai222d1 U2250 ( .A1(n7503), .A2(n784), .B1(n12575), .B2(n771), .C1(n7371), 
        .C2(1'b1), .ZN(n13642) );
  oai222d1 U2249 ( .A1(n7497), .A2(n784), .B1(n12574), .B2(n771), .C1(n7365), 
        .C2(1'b1), .ZN(n13641) );
  oai222d1 U2027 ( .A1(n7558), .A2(1'b1), .B1(n12372), .B2(n530), .C1(n7408), 
        .C2(n844), .ZN(n13439) );
  oai222d1 U2026 ( .A1(n7514), .A2(1'b1), .B1(n12371), .B2(n530), .C1(n7377), 
        .C2(n844), .ZN(n13438) );
  oai222d1 U2025 ( .A1(n7448), .A2(1'b1), .B1(n12370), .B2(n530), .C1(n7318), 
        .C2(n844), .ZN(n13437) );
  oai222d1 U2024 ( .A1(n7438), .A2(1'b1), .B1(n12369), .B2(n530), .C1(n7297), 
        .C2(n844), .ZN(n13436) );
  oai222d1 U2023 ( .A1(n7432), .A2(1'b1), .B1(n12368), .B2(n530), .C1(n7293), 
        .C2(n844), .ZN(n13435) );
  oai222d1 U2022 ( .A1(n7425), .A2(1'b1), .B1(n12367), .B2(n530), .C1(n7288), 
        .C2(n843), .ZN(n13434) );
  oai222d1 U2021 ( .A1(n7424), .A2(1'b1), .B1(n12366), .B2(n530), .C1(n7278), 
        .C2(n843), .ZN(n13433) );
  oai222d1 U2020 ( .A1(n7415), .A2(1'b1), .B1(n12365), .B2(n530), .C1(n7271), 
        .C2(n843), .ZN(n13432) );
  oai222d1 U2019 ( .A1(n7414), .A2(1'b1), .B1(n12364), .B2(n530), .C1(n7265), 
        .C2(n843), .ZN(n13431) );
  oai222d1 U2018 ( .A1(n7412), .A2(1'b1), .B1(n12363), .B2(n531), .C1(n7261), 
        .C2(n843), .ZN(n13430) );
  oai222d1 U2017 ( .A1(n7553), .A2(1'b1), .B1(n12362), .B2(n531), .C1(n7405), 
        .C2(n843), .ZN(n13429) );
  oai222d1 U2016 ( .A1(n7552), .A2(1'b1), .B1(n12361), .B2(n531), .C1(n7403), 
        .C2(n843), .ZN(n13428) );
  oai222d1 U2015 ( .A1(n7549), .A2(1'b1), .B1(n12360), .B2(n531), .C1(n7402), 
        .C2(n843), .ZN(n13427) );
  oai222d1 U2014 ( .A1(n7542), .A2(1'b1), .B1(n12359), .B2(n531), .C1(n7399), 
        .C2(n843), .ZN(n13426) );
  oai222d1 U2013 ( .A1(n7538), .A2(1'b1), .B1(n12358), .B2(n531), .C1(n7398), 
        .C2(n842), .ZN(n13425) );
  oai222d1 U2012 ( .A1(n7531), .A2(1'b1), .B1(n12357), .B2(n531), .C1(n7397), 
        .C2(n842), .ZN(n13424) );
  oai222d1 U2011 ( .A1(n7525), .A2(1'b1), .B1(n12356), .B2(n531), .C1(n7390), 
        .C2(n842), .ZN(n13423) );
  oai222d1 U2010 ( .A1(n7524), .A2(1'b1), .B1(n12355), .B2(n531), .C1(n7387), 
        .C2(n842), .ZN(n13422) );
  oai222d1 U2009 ( .A1(n7520), .A2(1'b1), .B1(n12354), .B2(n532), .C1(n7380), 
        .C2(n842), .ZN(n13421) );
  oai222d1 U2008 ( .A1(n7519), .A2(1'b1), .B1(n12353), .B2(n532), .C1(n7379), 
        .C2(n842), .ZN(n13420) );
  oai222d1 U2007 ( .A1(n7510), .A2(1'b1), .B1(n12352), .B2(n532), .C1(n7372), 
        .C2(n842), .ZN(n13419) );
  oai222d1 U2006 ( .A1(n7503), .A2(1'b1), .B1(n12351), .B2(n532), .C1(n7371), 
        .C2(n842), .ZN(n13418) );
  oai222d1 U2005 ( .A1(n7497), .A2(1'b1), .B1(n12350), .B2(n532), .C1(n7365), 
        .C2(n842), .ZN(n13417) );
  oai222d1 U2004 ( .A1(n7482), .A2(1'b1), .B1(n12349), .B2(n532), .C1(n7363), 
        .C2(n841), .ZN(n13416) );
  oai222d1 U2003 ( .A1(n7476), .A2(1'b1), .B1(n12348), .B2(n532), .C1(n7361), 
        .C2(n841), .ZN(n13415) );
  oai222d1 U2002 ( .A1(n7470), .A2(1'b1), .B1(n12347), .B2(n532), .C1(n7355), 
        .C2(n841), .ZN(n13414) );
  oai222d1 U2001 ( .A1(n7467), .A2(1'b1), .B1(n12346), .B2(n532), .C1(n7348), 
        .C2(n841), .ZN(n13413) );
  oai222d1 U2000 ( .A1(n7465), .A2(1'b1), .B1(n12345), .B2(n533), .C1(n7342), 
        .C2(n841), .ZN(n13412) );
  oai222d1 U1999 ( .A1(n7451), .A2(1'b1), .B1(n12344), .B2(n533), .C1(n7325), 
        .C2(n841), .ZN(n13411) );
  oai222d1 U1998 ( .A1(n7449), .A2(1'b1), .B1(n12343), .B2(n533), .C1(n7322), 
        .C2(n841), .ZN(n13410) );
  oai222d1 U1997 ( .A1(n7445), .A2(1'b1), .B1(n12342), .B2(n533), .C1(n7312), 
        .C2(n841), .ZN(n13409) );
  oai222d1 U1996 ( .A1(n7441), .A2(1'b1), .B1(n12341), .B2(n533), .C1(n7307), 
        .C2(n841), .ZN(n13408) );
  oai222d1 U1992 ( .A1(n7558), .A2(n861), .B1(n12340), .B2(n534), .C1(n7408), 
        .C2(1'b1), .ZN(n13407) );
  oai222d1 U1991 ( .A1(n7514), .A2(n861), .B1(n12339), .B2(n534), .C1(n7377), 
        .C2(1'b1), .ZN(n13406) );
  oai222d1 U1990 ( .A1(n7448), .A2(n861), .B1(n12338), .B2(n534), .C1(n7318), 
        .C2(1'b1), .ZN(n13405) );
  oai222d1 U1989 ( .A1(n7438), .A2(n861), .B1(n12337), .B2(n534), .C1(n7297), 
        .C2(1'b1), .ZN(n13404) );
  oai222d1 U1988 ( .A1(n7432), .A2(n861), .B1(n12336), .B2(n534), .C1(n7293), 
        .C2(1'b1), .ZN(n13403) );
  oai222d1 U1987 ( .A1(n7425), .A2(n861), .B1(n12335), .B2(n534), .C1(n7288), 
        .C2(1'b1), .ZN(n13402) );
  oai222d1 U1986 ( .A1(n7424), .A2(n861), .B1(n12334), .B2(n534), .C1(n7278), 
        .C2(1'b1), .ZN(n13401) );
  oai222d1 U1985 ( .A1(n7415), .A2(n861), .B1(n12333), .B2(n534), .C1(n7271), 
        .C2(1'b1), .ZN(n13400) );
  oai222d1 U1984 ( .A1(n7414), .A2(n860), .B1(n12332), .B2(n534), .C1(n7265), 
        .C2(1'b1), .ZN(n13399) );
  oai222d1 U1983 ( .A1(n7412), .A2(n860), .B1(n12331), .B2(n535), .C1(n7261), 
        .C2(1'b1), .ZN(n13398) );
  oai222d1 U1982 ( .A1(n7553), .A2(n860), .B1(n12330), .B2(n535), .C1(n7405), 
        .C2(1'b1), .ZN(n13397) );
  oai222d1 U1981 ( .A1(n7552), .A2(n860), .B1(n12329), .B2(n535), .C1(n7403), 
        .C2(1'b1), .ZN(n13396) );
  oai222d1 U1980 ( .A1(n7549), .A2(n860), .B1(n12328), .B2(n535), .C1(n7402), 
        .C2(1'b1), .ZN(n13395) );
  oai222d1 U1979 ( .A1(n7542), .A2(n860), .B1(n12327), .B2(n535), .C1(n7399), 
        .C2(1'b1), .ZN(n13394) );
  oai222d1 U1978 ( .A1(n7538), .A2(n860), .B1(n12326), .B2(n535), .C1(n7398), 
        .C2(1'b1), .ZN(n13393) );
  oai222d1 U1977 ( .A1(n7531), .A2(n860), .B1(n12325), .B2(n535), .C1(n7397), 
        .C2(1'b1), .ZN(n13392) );
  oai222d1 U1976 ( .A1(n7525), .A2(n860), .B1(n12324), .B2(n535), .C1(n7390), 
        .C2(1'b1), .ZN(n13391) );
  oai222d1 U1975 ( .A1(n7524), .A2(n860), .B1(n12323), .B2(n535), .C1(n7387), 
        .C2(1'b1), .ZN(n13390) );
  oai222d1 U1974 ( .A1(n7520), .A2(n859), .B1(n12322), .B2(n536), .C1(n7380), 
        .C2(1'b1), .ZN(n13389) );
  oai222d1 U1973 ( .A1(n7519), .A2(n859), .B1(n12321), .B2(n536), .C1(n7379), 
        .C2(1'b1), .ZN(n13388) );
  oai222d1 U1972 ( .A1(n7510), .A2(n859), .B1(n12320), .B2(n536), .C1(n7372), 
        .C2(1'b1), .ZN(n13387) );
  oai222d1 U1971 ( .A1(n7503), .A2(n859), .B1(n12319), .B2(n536), .C1(n7371), 
        .C2(1'b1), .ZN(n13386) );
  oai222d1 U1970 ( .A1(n7497), .A2(n859), .B1(n12318), .B2(n536), .C1(n7365), 
        .C2(1'b1), .ZN(n13385) );
  oai222d1 U1969 ( .A1(n7482), .A2(n859), .B1(n12317), .B2(n536), .C1(n7363), 
        .C2(1'b1), .ZN(n13384) );
  oai222d1 U1968 ( .A1(n7476), .A2(n859), .B1(n12316), .B2(n536), .C1(n7361), 
        .C2(1'b1), .ZN(n13383) );
  oai222d1 U1967 ( .A1(n7470), .A2(n859), .B1(n12315), .B2(n536), .C1(n7355), 
        .C2(1'b1), .ZN(n13382) );
  oai222d1 U1966 ( .A1(n7467), .A2(n859), .B1(n12314), .B2(n536), .C1(n7348), 
        .C2(1'b1), .ZN(n13381) );
  oai222d1 U1965 ( .A1(n7465), .A2(n859), .B1(n12313), .B2(n537), .C1(n7342), 
        .C2(1'b1), .ZN(n13380) );
  oai222d1 U1964 ( .A1(n7451), .A2(n858), .B1(n12312), .B2(n537), .C1(n7325), 
        .C2(1'b1), .ZN(n13379) );
  oai222d1 U1963 ( .A1(n7449), .A2(n858), .B1(n12311), .B2(n537), .C1(n7322), 
        .C2(1'b1), .ZN(n13378) );
  oai222d1 U1962 ( .A1(n7445), .A2(n858), .B1(n12310), .B2(n537), .C1(n7312), 
        .C2(1'b1), .ZN(n13377) );
  oai222d1 U1961 ( .A1(n7441), .A2(n858), .B1(n12309), .B2(n537), .C1(n7307), 
        .C2(1'b1), .ZN(n13376) );
  oai222d1 U2248 ( .A1(n7482), .A2(n784), .B1(n12573), .B2(n771), .C1(n7363), 
        .C2(1'b1), .ZN(n13640) );
  oai222d1 U2247 ( .A1(n7476), .A2(n784), .B1(n12572), .B2(n771), .C1(n7361), 
        .C2(1'b1), .ZN(n13639) );
  oai222d1 U2246 ( .A1(n7470), .A2(n784), .B1(n12571), .B2(n771), .C1(n7355), 
        .C2(1'b1), .ZN(n13638) );
  oai222d1 U2245 ( .A1(n7467), .A2(n784), .B1(n12570), .B2(n771), .C1(n7348), 
        .C2(1'b1), .ZN(n13637) );
  oai222d1 U2244 ( .A1(n7465), .A2(n785), .B1(n12569), .B2(n772), .C1(n7342), 
        .C2(1'b1), .ZN(n13636) );
  oai222d1 U2243 ( .A1(n7451), .A2(n785), .B1(n12568), .B2(n772), .C1(n7325), 
        .C2(1'b1), .ZN(n13635) );
  oai222d1 U2242 ( .A1(n7449), .A2(n785), .B1(n12567), .B2(n772), .C1(n7322), 
        .C2(1'b1), .ZN(n13634) );
  oai222d1 U2241 ( .A1(n7445), .A2(n785), .B1(n12566), .B2(n772), .C1(n7312), 
        .C2(1'b1), .ZN(n13633) );
  oai222d1 U2240 ( .A1(n7441), .A2(n785), .B1(n12565), .B2(n772), .C1(n7307), 
        .C2(1'b1), .ZN(n13632) );
  oai222d1 U2176 ( .A1(n7441), .A2(n806), .B1(n12501), .B2(n802), .C1(n7307), 
        .C2(1'b1), .ZN(n13569) );
  oai222d1 U2376 ( .A1(n7558), .A2(1'b1), .B1(n12692), .B2(n727), .C1(n7408), 
        .C2(n721), .ZN(n13759) );
  oai222d1 U2375 ( .A1(n7514), .A2(1'b1), .B1(n12691), .B2(n727), .C1(n7377), 
        .C2(n721), .ZN(n13758) );
  oai222d1 U2374 ( .A1(n7448), .A2(1'b1), .B1(n12690), .B2(n727), .C1(n7318), 
        .C2(n721), .ZN(n13757) );
  oai222d1 U2373 ( .A1(n7438), .A2(1'b1), .B1(n12689), .B2(n727), .C1(n7297), 
        .C2(n721), .ZN(n13756) );
  oai222d1 U2372 ( .A1(n7432), .A2(1'b1), .B1(n12688), .B2(n727), .C1(n7293), 
        .C2(n721), .ZN(n13755) );
  oai222d1 U2371 ( .A1(n7425), .A2(1'b1), .B1(n12687), .B2(n727), .C1(n7288), 
        .C2(n720), .ZN(n13754) );
  oai222d1 U2370 ( .A1(n7424), .A2(1'b1), .B1(n12686), .B2(n727), .C1(n7278), 
        .C2(n720), .ZN(n13753) );
  oai222d1 U2369 ( .A1(n7415), .A2(1'b1), .B1(n12685), .B2(n727), .C1(n7271), 
        .C2(n720), .ZN(n13752) );
  oai222d1 U2368 ( .A1(n7414), .A2(1'b1), .B1(n12684), .B2(n727), .C1(n7265), 
        .C2(n720), .ZN(n13751) );
  oai222d1 U2367 ( .A1(n7412), .A2(1'b1), .B1(n12683), .B2(n728), .C1(n7261), 
        .C2(n720), .ZN(n13750) );
  oai222d1 U2366 ( .A1(n7553), .A2(1'b1), .B1(n12682), .B2(n728), .C1(n7405), 
        .C2(n720), .ZN(n13749) );
  oai222d1 U2365 ( .A1(n7552), .A2(1'b1), .B1(n12681), .B2(n728), .C1(n7403), 
        .C2(n720), .ZN(n13748) );
  oai222d1 U2364 ( .A1(n7549), .A2(1'b1), .B1(n12680), .B2(n728), .C1(n7402), 
        .C2(n720), .ZN(n13747) );
  oai222d1 U2363 ( .A1(n7542), .A2(1'b1), .B1(n12679), .B2(n728), .C1(n7399), 
        .C2(n720), .ZN(n13746) );
  oai222d1 U2362 ( .A1(n7538), .A2(1'b1), .B1(n12678), .B2(n728), .C1(n7398), 
        .C2(n719), .ZN(n13745) );
  oai222d1 U2361 ( .A1(n7531), .A2(1'b1), .B1(n12677), .B2(n728), .C1(n7397), 
        .C2(n719), .ZN(n13744) );
  oai222d1 U2360 ( .A1(n7525), .A2(1'b1), .B1(n12676), .B2(n728), .C1(n7390), 
        .C2(n719), .ZN(n13743) );
  oai222d1 U2359 ( .A1(n7524), .A2(1'b1), .B1(n12675), .B2(n728), .C1(n7387), 
        .C2(n719), .ZN(n13742) );
  oai222d1 U2358 ( .A1(n7520), .A2(1'b1), .B1(n12674), .B2(n729), .C1(n7380), 
        .C2(n719), .ZN(n13741) );
  oai222d1 U2357 ( .A1(n7519), .A2(1'b1), .B1(n12673), .B2(n729), .C1(n7379), 
        .C2(n719), .ZN(n13740) );
  oai222d1 U2356 ( .A1(n7510), .A2(1'b1), .B1(n12672), .B2(n729), .C1(n7372), 
        .C2(n719), .ZN(n13739) );
  oai222d1 U2355 ( .A1(n7503), .A2(1'b1), .B1(n12671), .B2(n729), .C1(n7371), 
        .C2(n719), .ZN(n13738) );
  oai222d1 U2354 ( .A1(n7497), .A2(1'b1), .B1(n12670), .B2(n729), .C1(n7365), 
        .C2(n719), .ZN(n13737) );
  oai222d1 U2353 ( .A1(n7482), .A2(1'b1), .B1(n12669), .B2(n729), .C1(n7363), 
        .C2(n718), .ZN(n13736) );
  oai222d1 U2352 ( .A1(n7476), .A2(1'b1), .B1(n12668), .B2(n729), .C1(n7361), 
        .C2(n718), .ZN(n13735) );
  oai222d1 U2351 ( .A1(n7470), .A2(1'b1), .B1(n12667), .B2(n729), .C1(n7355), 
        .C2(n718), .ZN(n13734) );
  oai222d1 U2350 ( .A1(n7467), .A2(1'b1), .B1(n12666), .B2(n729), .C1(n7348), 
        .C2(n718), .ZN(n13733) );
  oai222d1 U2349 ( .A1(n7465), .A2(1'b1), .B1(n12665), .B2(n730), .C1(n7342), 
        .C2(n718), .ZN(n13732) );
  oai222d1 U2348 ( .A1(n7451), .A2(1'b1), .B1(n12664), .B2(n730), .C1(n7325), 
        .C2(n718), .ZN(n13731) );
  oai222d1 U2347 ( .A1(n7449), .A2(1'b1), .B1(n12663), .B2(n730), .C1(n7322), 
        .C2(n718), .ZN(n13730) );
  oai222d1 U2346 ( .A1(n7445), .A2(1'b1), .B1(n12662), .B2(n730), .C1(n7312), 
        .C2(n718), .ZN(n13729) );
  oai222d1 U2345 ( .A1(n7441), .A2(1'b1), .B1(n12661), .B2(n730), .C1(n7307), 
        .C2(n718), .ZN(n13728) );
  oai222d1 U2341 ( .A1(n7558), .A2(n753), .B1(n12660), .B2(n740), .C1(n7408), 
        .C2(1'b1), .ZN(n13727) );
  oai222d1 U2340 ( .A1(n7514), .A2(n753), .B1(n12659), .B2(n740), .C1(n7377), 
        .C2(1'b1), .ZN(n13726) );
  oai222d1 U2339 ( .A1(n7448), .A2(n753), .B1(n12658), .B2(n740), .C1(n7318), 
        .C2(1'b1), .ZN(n13725) );
  oai222d1 U2338 ( .A1(n7438), .A2(n753), .B1(n12657), .B2(n740), .C1(n7297), 
        .C2(1'b1), .ZN(n13724) );
  oai222d1 U2337 ( .A1(n7432), .A2(n753), .B1(n12656), .B2(n740), .C1(n7293), 
        .C2(1'b1), .ZN(n13723) );
  oai222d1 U2336 ( .A1(n7425), .A2(n753), .B1(n12655), .B2(n740), .C1(n7288), 
        .C2(1'b1), .ZN(n13722) );
  oai222d1 U2335 ( .A1(n7424), .A2(n753), .B1(n12654), .B2(n740), .C1(n7278), 
        .C2(1'b1), .ZN(n13721) );
  oai222d1 U2334 ( .A1(n7415), .A2(n753), .B1(n12653), .B2(n740), .C1(n7271), 
        .C2(1'b1), .ZN(n13720) );
  oai222d1 U2333 ( .A1(n7414), .A2(n752), .B1(n12652), .B2(n740), .C1(n7265), 
        .C2(1'b1), .ZN(n13719) );
  oai222d1 U2332 ( .A1(n7412), .A2(n752), .B1(n12651), .B2(n741), .C1(n7261), 
        .C2(1'b1), .ZN(n13718) );
  oai222d1 U2331 ( .A1(n7553), .A2(n752), .B1(n12650), .B2(n741), .C1(n7405), 
        .C2(1'b1), .ZN(n13717) );
  oai222d1 U2330 ( .A1(n7552), .A2(n752), .B1(n12649), .B2(n741), .C1(n7403), 
        .C2(1'b1), .ZN(n13716) );
  oai222d1 U2329 ( .A1(n7549), .A2(n752), .B1(n12648), .B2(n741), .C1(n7402), 
        .C2(1'b1), .ZN(n13715) );
  oai222d1 U2328 ( .A1(n7542), .A2(n752), .B1(n12647), .B2(n741), .C1(n7399), 
        .C2(1'b1), .ZN(n13714) );
  oai222d1 U2327 ( .A1(n7538), .A2(n752), .B1(n12646), .B2(n741), .C1(n7398), 
        .C2(1'b1), .ZN(n13713) );
  oai222d1 U2326 ( .A1(n7531), .A2(n752), .B1(n12645), .B2(n741), .C1(n7397), 
        .C2(1'b1), .ZN(n13712) );
  oai222d1 U2325 ( .A1(n7525), .A2(n752), .B1(n12644), .B2(n741), .C1(n7390), 
        .C2(1'b1), .ZN(n13711) );
  oai222d1 U2324 ( .A1(n7524), .A2(n752), .B1(n12643), .B2(n741), .C1(n7387), 
        .C2(1'b1), .ZN(n13710) );
  oai222d1 U2323 ( .A1(n7520), .A2(n751), .B1(n12642), .B2(n742), .C1(n7380), 
        .C2(1'b1), .ZN(n13709) );
  oai222d1 U2322 ( .A1(n7519), .A2(n751), .B1(n12641), .B2(n742), .C1(n7379), 
        .C2(1'b1), .ZN(n13708) );
  oai222d1 U2321 ( .A1(n7510), .A2(n751), .B1(n12640), .B2(n742), .C1(n7372), 
        .C2(1'b1), .ZN(n13707) );
  oai222d1 U2320 ( .A1(n7503), .A2(n751), .B1(n12639), .B2(n742), .C1(n7371), 
        .C2(1'b1), .ZN(n13706) );
  oai222d1 U2319 ( .A1(n7497), .A2(n751), .B1(n12638), .B2(n742), .C1(n7365), 
        .C2(1'b1), .ZN(n13705) );
  oai222d1 U2097 ( .A1(n7558), .A2(1'b1), .B1(n12436), .B2(n522), .C1(n7408), 
        .C2(n827), .ZN(n13503) );
  oai222d1 U2096 ( .A1(n7514), .A2(1'b1), .B1(n12435), .B2(n522), .C1(n7377), 
        .C2(n827), .ZN(n13502) );
  oai222d1 U2095 ( .A1(n7448), .A2(1'b1), .B1(n12434), .B2(n522), .C1(n7318), 
        .C2(n827), .ZN(n13501) );
  oai222d1 U2094 ( .A1(n7438), .A2(1'b1), .B1(n12433), .B2(n522), .C1(n7297), 
        .C2(n827), .ZN(n13500) );
  oai222d1 U2093 ( .A1(n7432), .A2(1'b1), .B1(n12432), .B2(n522), .C1(n7293), 
        .C2(n827), .ZN(n13499) );
  oai222d1 U2092 ( .A1(n7425), .A2(1'b1), .B1(n12431), .B2(n522), .C1(n7288), 
        .C2(n826), .ZN(n13498) );
  oai222d1 U2091 ( .A1(n7424), .A2(1'b1), .B1(n12430), .B2(n522), .C1(n7278), 
        .C2(n826), .ZN(n13497) );
  oai222d1 U2090 ( .A1(n7415), .A2(1'b1), .B1(n12429), .B2(n522), .C1(n7271), 
        .C2(n826), .ZN(n13496) );
  oai222d1 U2089 ( .A1(n7414), .A2(1'b1), .B1(n12428), .B2(n522), .C1(n7265), 
        .C2(n826), .ZN(n13495) );
  oai222d1 U2088 ( .A1(n7412), .A2(1'b1), .B1(n12427), .B2(n523), .C1(n7261), 
        .C2(n826), .ZN(n13494) );
  oai222d1 U2087 ( .A1(n7553), .A2(1'b1), .B1(n12426), .B2(n523), .C1(n7405), 
        .C2(n826), .ZN(n13493) );
  oai222d1 U2086 ( .A1(n7552), .A2(1'b1), .B1(n12425), .B2(n523), .C1(n7403), 
        .C2(n826), .ZN(n13492) );
  oai222d1 U2085 ( .A1(n7549), .A2(1'b1), .B1(n12424), .B2(n523), .C1(n7402), 
        .C2(n826), .ZN(n13491) );
  oai222d1 U2084 ( .A1(n7542), .A2(1'b1), .B1(n12423), .B2(n523), .C1(n7399), 
        .C2(n826), .ZN(n13490) );
  oai222d1 U2083 ( .A1(n7538), .A2(1'b1), .B1(n12422), .B2(n523), .C1(n7398), 
        .C2(n825), .ZN(n13489) );
  oai222d1 U2082 ( .A1(n7531), .A2(1'b1), .B1(n12421), .B2(n523), .C1(n7397), 
        .C2(n825), .ZN(n13488) );
  oai222d1 U2081 ( .A1(n7525), .A2(1'b1), .B1(n12420), .B2(n523), .C1(n7390), 
        .C2(n825), .ZN(n13487) );
  oai222d1 U2080 ( .A1(n7524), .A2(1'b1), .B1(n12419), .B2(n523), .C1(n7387), 
        .C2(n825), .ZN(n13486) );
  oai222d1 U2079 ( .A1(n7520), .A2(1'b1), .B1(n12418), .B2(n524), .C1(n7380), 
        .C2(n825), .ZN(n13485) );
  oai222d1 U2078 ( .A1(n7519), .A2(1'b1), .B1(n12417), .B2(n524), .C1(n7379), 
        .C2(n825), .ZN(n13484) );
  oai222d1 U2077 ( .A1(n7510), .A2(1'b1), .B1(n12416), .B2(n524), .C1(n7372), 
        .C2(n825), .ZN(n13483) );
  oai222d1 U2076 ( .A1(n7503), .A2(1'b1), .B1(n12415), .B2(n524), .C1(n7371), 
        .C2(n825), .ZN(n13482) );
  oai222d1 U2075 ( .A1(n7497), .A2(1'b1), .B1(n12414), .B2(n524), .C1(n7365), 
        .C2(n825), .ZN(n13481) );
  oai222d1 U2074 ( .A1(n7482), .A2(1'b1), .B1(n12413), .B2(n524), .C1(n7363), 
        .C2(n824), .ZN(n13480) );
  oai222d1 U2073 ( .A1(n7476), .A2(1'b1), .B1(n12412), .B2(n524), .C1(n7361), 
        .C2(n824), .ZN(n13479) );
  oai222d1 U2072 ( .A1(n7470), .A2(1'b1), .B1(n12411), .B2(n524), .C1(n7355), 
        .C2(n824), .ZN(n13478) );
  oai222d1 U2071 ( .A1(n7467), .A2(1'b1), .B1(n12410), .B2(n524), .C1(n7348), 
        .C2(n824), .ZN(n13477) );
  oai222d1 U2070 ( .A1(n7465), .A2(1'b1), .B1(n12409), .B2(n525), .C1(n7342), 
        .C2(n824), .ZN(n13476) );
  oai222d1 U2069 ( .A1(n7451), .A2(1'b1), .B1(n12408), .B2(n525), .C1(n7325), 
        .C2(n824), .ZN(n13475) );
  oai222d1 U2068 ( .A1(n7449), .A2(1'b1), .B1(n12407), .B2(n525), .C1(n7322), 
        .C2(n824), .ZN(n13474) );
  oai222d1 U2067 ( .A1(n7445), .A2(1'b1), .B1(n12406), .B2(n525), .C1(n7312), 
        .C2(n824), .ZN(n13473) );
  oai222d1 U2066 ( .A1(n7441), .A2(1'b1), .B1(n12405), .B2(n525), .C1(n7307), 
        .C2(n824), .ZN(n13472) );
  oai222d1 U2062 ( .A1(n7558), .A2(n847), .B1(n12404), .B2(n526), .C1(n7408), 
        .C2(1'b1), .ZN(n13471) );
  oai222d1 U2061 ( .A1(n7514), .A2(n847), .B1(n12403), .B2(n526), .C1(n7377), 
        .C2(1'b1), .ZN(n13470) );
  oai222d1 U2060 ( .A1(n7448), .A2(n847), .B1(n12402), .B2(n526), .C1(n7318), 
        .C2(1'b1), .ZN(n13469) );
  oai222d1 U2059 ( .A1(n7438), .A2(n847), .B1(n12401), .B2(n526), .C1(n7297), 
        .C2(1'b1), .ZN(n13468) );
  oai222d1 U2058 ( .A1(n7432), .A2(n847), .B1(n12400), .B2(n526), .C1(n7293), 
        .C2(1'b1), .ZN(n13467) );
  oai222d1 U2057 ( .A1(n7425), .A2(n847), .B1(n12399), .B2(n526), .C1(n7288), 
        .C2(1'b1), .ZN(n13466) );
  oai222d1 U2056 ( .A1(n7424), .A2(n847), .B1(n12398), .B2(n526), .C1(n7278), 
        .C2(1'b1), .ZN(n13465) );
  oai222d1 U2055 ( .A1(n7415), .A2(n847), .B1(n12397), .B2(n526), .C1(n7271), 
        .C2(1'b1), .ZN(n13464) );
  oai222d1 U2054 ( .A1(n7414), .A2(n846), .B1(n12396), .B2(n526), .C1(n7265), 
        .C2(1'b1), .ZN(n13463) );
  oai222d1 U2053 ( .A1(n7412), .A2(n846), .B1(n12395), .B2(n527), .C1(n7261), 
        .C2(1'b1), .ZN(n13462) );
  oai222d1 U2052 ( .A1(n7553), .A2(n846), .B1(n12394), .B2(n527), .C1(n7405), 
        .C2(1'b1), .ZN(n13461) );
  oai222d1 U2051 ( .A1(n7552), .A2(n846), .B1(n12393), .B2(n527), .C1(n7403), 
        .C2(1'b1), .ZN(n13460) );
  oai222d1 U2050 ( .A1(n7549), .A2(n846), .B1(n12392), .B2(n527), .C1(n7402), 
        .C2(1'b1), .ZN(n13459) );
  oai222d1 U2049 ( .A1(n7542), .A2(n846), .B1(n12391), .B2(n527), .C1(n7399), 
        .C2(1'b1), .ZN(n13458) );
  oai222d1 U2048 ( .A1(n7538), .A2(n846), .B1(n12390), .B2(n527), .C1(n7398), 
        .C2(1'b1), .ZN(n13457) );
  oai222d1 U2047 ( .A1(n7531), .A2(n846), .B1(n12389), .B2(n527), .C1(n7397), 
        .C2(1'b1), .ZN(n13456) );
  oai222d1 U2046 ( .A1(n7525), .A2(n846), .B1(n12388), .B2(n527), .C1(n7390), 
        .C2(1'b1), .ZN(n13455) );
  oai222d1 U2045 ( .A1(n7524), .A2(n846), .B1(n12387), .B2(n527), .C1(n7387), 
        .C2(1'b1), .ZN(n13454) );
  oai222d1 U2044 ( .A1(n7520), .A2(n845), .B1(n12386), .B2(n528), .C1(n7380), 
        .C2(1'b1), .ZN(n13453) );
  oai222d1 U2043 ( .A1(n7519), .A2(n845), .B1(n12385), .B2(n528), .C1(n7379), 
        .C2(1'b1), .ZN(n13452) );
  oai222d1 U2042 ( .A1(n7510), .A2(n845), .B1(n12384), .B2(n528), .C1(n7372), 
        .C2(1'b1), .ZN(n13451) );
  oai222d1 U2041 ( .A1(n7503), .A2(n845), .B1(n12383), .B2(n528), .C1(n7371), 
        .C2(1'b1), .ZN(n13450) );
  oai222d1 U2040 ( .A1(n7497), .A2(n845), .B1(n12382), .B2(n528), .C1(n7365), 
        .C2(1'b1), .ZN(n13449) );
  oai222d1 U2039 ( .A1(n7482), .A2(n845), .B1(n12381), .B2(n528), .C1(n7363), 
        .C2(1'b1), .ZN(n13448) );
  oai222d1 U2038 ( .A1(n7476), .A2(n845), .B1(n12380), .B2(n528), .C1(n7361), 
        .C2(1'b1), .ZN(n13447) );
  oai222d1 U2037 ( .A1(n7470), .A2(n845), .B1(n12379), .B2(n528), .C1(n7355), 
        .C2(1'b1), .ZN(n13446) );
  oai222d1 U2036 ( .A1(n7467), .A2(n845), .B1(n12378), .B2(n528), .C1(n7348), 
        .C2(1'b1), .ZN(n13445) );
  oai222d1 U2035 ( .A1(n7465), .A2(n845), .B1(n12377), .B2(n529), .C1(n7342), 
        .C2(1'b1), .ZN(n13444) );
  oai222d1 U2034 ( .A1(n7451), .A2(n844), .B1(n12376), .B2(n529), .C1(n7325), 
        .C2(1'b1), .ZN(n13443) );
  oai222d1 U2033 ( .A1(n7449), .A2(n844), .B1(n12375), .B2(n529), .C1(n7322), 
        .C2(1'b1), .ZN(n13442) );
  oai222d1 U2032 ( .A1(n7445), .A2(n844), .B1(n12374), .B2(n529), .C1(n7312), 
        .C2(1'b1), .ZN(n13441) );
  oai222d1 U2031 ( .A1(n7441), .A2(n844), .B1(n12373), .B2(n529), .C1(n7307), 
        .C2(1'b1), .ZN(n13440) );
  oai222d1 U2318 ( .A1(n7482), .A2(n751), .B1(n12637), .B2(n742), .C1(n7363), 
        .C2(1'b1), .ZN(n13704) );
  oai222d1 U2317 ( .A1(n7476), .A2(n751), .B1(n12636), .B2(n742), .C1(n7361), 
        .C2(1'b1), .ZN(n13703) );
  oai222d1 U2316 ( .A1(n7470), .A2(n751), .B1(n12635), .B2(n742), .C1(n7355), 
        .C2(1'b1), .ZN(n13702) );
  oai222d1 U2315 ( .A1(n7467), .A2(n751), .B1(n12634), .B2(n742), .C1(n7348), 
        .C2(1'b1), .ZN(n13701) );
  oai222d1 U2314 ( .A1(n7465), .A2(n751), .B1(n12633), .B2(n743), .C1(n7342), 
        .C2(1'b1), .ZN(n13700) );
  oai222d1 U2313 ( .A1(n7451), .A2(n750), .B1(n12632), .B2(n743), .C1(n7325), 
        .C2(1'b1), .ZN(n13699) );
  oai222d1 U2312 ( .A1(n7449), .A2(n750), .B1(n12631), .B2(n743), .C1(n7322), 
        .C2(1'b1), .ZN(n13698) );
  oai222d1 U2311 ( .A1(n7445), .A2(n750), .B1(n12630), .B2(n743), .C1(n7312), 
        .C2(1'b1), .ZN(n13697) );
  oai222d1 U2310 ( .A1(n7441), .A2(n750), .B1(n12629), .B2(n743), .C1(n7307), 
        .C2(1'b1), .ZN(n13696) );
  oai222d1 U2177 ( .A1(n7445), .A2(n806), .B1(n12502), .B2(n802), .C1(n7312), 
        .C2(1'b1), .ZN(n13570) );
  oai222d1 U2178 ( .A1(n7449), .A2(n806), .B1(n12503), .B2(n802), .C1(n7322), 
        .C2(1'b1), .ZN(n13571) );
  oai222d1 U2179 ( .A1(n7451), .A2(n806), .B1(n12504), .B2(n802), .C1(n7325), 
        .C2(1'b1), .ZN(n13572) );
  oai222d1 U2180 ( .A1(n7465), .A2(n807), .B1(n12505), .B2(n802), .C1(n7342), 
        .C2(1'b1), .ZN(n13573) );
  oai222d1 U2181 ( .A1(n7467), .A2(n807), .B1(n12506), .B2(n801), .C1(n7348), 
        .C2(1'b1), .ZN(n13574) );
  oai222d1 U2182 ( .A1(n7470), .A2(n807), .B1(n12507), .B2(n801), .C1(n7355), 
        .C2(1'b1), .ZN(n13575) );
  oai222d1 U2183 ( .A1(n7476), .A2(n807), .B1(n12508), .B2(n801), .C1(n7361), 
        .C2(1'b1), .ZN(n13576) );
  oai222d1 U2184 ( .A1(n7482), .A2(n807), .B1(n12509), .B2(n801), .C1(n7363), 
        .C2(1'b1), .ZN(n13577) );
  oai222d1 U2185 ( .A1(n7497), .A2(n807), .B1(n12510), .B2(n801), .C1(n7365), 
        .C2(1'b1), .ZN(n13578) );
  oai222d1 U2186 ( .A1(n7503), .A2(n807), .B1(n12511), .B2(n801), .C1(n7371), 
        .C2(1'b1), .ZN(n13579) );
  oai222d1 U2187 ( .A1(n7510), .A2(n807), .B1(n12512), .B2(n801), .C1(n7372), 
        .C2(1'b1), .ZN(n13580) );
  oai222d1 U2188 ( .A1(n7519), .A2(n807), .B1(n12513), .B2(n801), .C1(n7379), 
        .C2(1'b1), .ZN(n13581) );
  oai222d1 U2189 ( .A1(n7520), .A2(n807), .B1(n12514), .B2(n801), .C1(n7380), 
        .C2(1'b1), .ZN(n13582) );
  oai222d1 U2190 ( .A1(n7524), .A2(n808), .B1(n12515), .B2(n800), .C1(n7387), 
        .C2(1'b1), .ZN(n13583) );
  oai222d1 U2191 ( .A1(n7525), .A2(n808), .B1(n12516), .B2(n800), .C1(n7390), 
        .C2(1'b1), .ZN(n13584) );
  oai222d1 U2192 ( .A1(n7531), .A2(n808), .B1(n12517), .B2(n800), .C1(n7397), 
        .C2(1'b1), .ZN(n13585) );
  oai222d1 U2193 ( .A1(n7538), .A2(n808), .B1(n12518), .B2(n800), .C1(n7398), 
        .C2(1'b1), .ZN(n13586) );
  oai222d1 U2194 ( .A1(n7542), .A2(n808), .B1(n12519), .B2(n800), .C1(n7399), 
        .C2(1'b1), .ZN(n13587) );
  oai222d1 U2195 ( .A1(n7549), .A2(n808), .B1(n12520), .B2(n800), .C1(n7402), 
        .C2(1'b1), .ZN(n13588) );
  oai222d1 U2196 ( .A1(n7552), .A2(n808), .B1(n12521), .B2(n800), .C1(n7403), 
        .C2(1'b1), .ZN(n13589) );
  oai222d1 U2197 ( .A1(n7553), .A2(n808), .B1(n12522), .B2(n800), .C1(n7405), 
        .C2(1'b1), .ZN(n13590) );
  oai222d1 U2198 ( .A1(n7412), .A2(n808), .B1(n12523), .B2(n800), .C1(n7261), 
        .C2(1'b1), .ZN(n13591) );
  oai222d1 U2199 ( .A1(n7414), .A2(n808), .B1(n12524), .B2(n799), .C1(n7265), 
        .C2(1'b1), .ZN(n13592) );
  oai222d1 U2200 ( .A1(n7415), .A2(n809), .B1(n12525), .B2(n799), .C1(n7271), 
        .C2(1'b1), .ZN(n13593) );
  oai222d1 U2201 ( .A1(n7424), .A2(n809), .B1(n12526), .B2(n799), .C1(n7278), 
        .C2(1'b1), .ZN(n13594) );
  oai222d1 U2202 ( .A1(n7425), .A2(n809), .B1(n12527), .B2(n799), .C1(n7288), 
        .C2(1'b1), .ZN(n13595) );
  oai222d1 U2203 ( .A1(n7438), .A2(n809), .B1(n12529), .B2(n799), .C1(n7297), 
        .C2(1'b1), .ZN(n13596) );
  oai222d1 U2204 ( .A1(n7448), .A2(n809), .B1(n12530), .B2(n799), .C1(n7318), 
        .C2(1'b1), .ZN(n13597) );
  oai222d1 U2205 ( .A1(n7514), .A2(n809), .B1(n12531), .B2(n799), .C1(n7377), 
        .C2(1'b1), .ZN(n13598) );
  oai222d1 U2206 ( .A1(n7558), .A2(n809), .B1(n12532), .B2(n799), .C1(n7408), 
        .C2(1'b1), .ZN(n13599) );
  oai222d1 U2207 ( .A1(n7307), .A2(n781), .B1(n12533), .B2(n778), .C1(n7441), 
        .C2(1'b1), .ZN(n13600) );
  oai222d1 U2208 ( .A1(n7312), .A2(n788), .B1(n12534), .B2(n778), .C1(n7445), 
        .C2(1'b1), .ZN(n13601) );
  oai222d1 U2209 ( .A1(n7322), .A2(n788), .B1(n12535), .B2(n778), .C1(n7449), 
        .C2(1'b1), .ZN(n13602) );
  oai222d1 U2210 ( .A1(n7325), .A2(n788), .B1(n12536), .B2(n778), .C1(n7451), 
        .C2(1'b1), .ZN(n13603) );
  oai222d1 U2211 ( .A1(n7342), .A2(n788), .B1(n12537), .B2(n778), .C1(n7465), 
        .C2(1'b1), .ZN(n13604) );
  oai222d1 U2212 ( .A1(n7348), .A2(n788), .B1(n12538), .B2(n777), .C1(n7467), 
        .C2(1'b1), .ZN(n13605) );
  oai222d1 U1947 ( .A1(n7553), .A2(1'b1), .B1(n12298), .B2(n539), .C1(n7405), 
        .C2(n857), .ZN(n13365) );
  oai222d1 U1946 ( .A1(n7552), .A2(1'b1), .B1(n12297), .B2(n539), .C1(n7403), 
        .C2(n857), .ZN(n13364) );
  oai222d1 U1951 ( .A1(n7424), .A2(1'b1), .B1(n12302), .B2(n538), .C1(n7278), 
        .C2(n857), .ZN(n13369) );
  oai222d1 U1944 ( .A1(n7542), .A2(1'b1), .B1(n12295), .B2(n539), .C1(n7399), 
        .C2(n857), .ZN(n13362) );
  oai222d1 U1943 ( .A1(n7538), .A2(1'b1), .B1(n12294), .B2(n539), .C1(n7398), 
        .C2(n856), .ZN(n13361) );
  oai222d1 U1942 ( .A1(n7531), .A2(1'b1), .B1(n12293), .B2(n539), .C1(n7397), 
        .C2(n856), .ZN(n13360) );
  oai222d1 U1941 ( .A1(n7525), .A2(1'b1), .B1(n12292), .B2(n539), .C1(n7390), 
        .C2(n856), .ZN(n13359) );
  oai222d1 U1940 ( .A1(n7524), .A2(1'b1), .B1(n12291), .B2(n539), .C1(n7387), 
        .C2(n856), .ZN(n13358) );
  oai222d1 U1945 ( .A1(n7549), .A2(1'b1), .B1(n12296), .B2(n539), .C1(n7402), 
        .C2(n857), .ZN(n13363) );
  oai222d1 U1938 ( .A1(n7519), .A2(1'b1), .B1(n12289), .B2(n540), .C1(n7379), 
        .C2(n856), .ZN(n13356) );
  oai222d1 U1937 ( .A1(n7510), .A2(1'b1), .B1(n12288), .B2(n540), .C1(n7372), 
        .C2(n856), .ZN(n13355) );
  oai222d1 U1936 ( .A1(n7503), .A2(1'b1), .B1(n12287), .B2(n540), .C1(n7371), 
        .C2(n856), .ZN(n13354) );
  oai222d1 U1935 ( .A1(n7497), .A2(1'b1), .B1(n12286), .B2(n540), .C1(n7365), 
        .C2(n856), .ZN(n13353) );
  oai222d1 U1934 ( .A1(n7482), .A2(1'b1), .B1(n12285), .B2(n540), .C1(n7363), 
        .C2(n855), .ZN(n13352) );
  oai222d1 U1939 ( .A1(n7520), .A2(1'b1), .B1(n12290), .B2(n540), .C1(n7380), 
        .C2(n856), .ZN(n13357) );
  oai222d1 U1932 ( .A1(n7470), .A2(1'b1), .B1(n12283), .B2(n540), .C1(n7355), 
        .C2(n855), .ZN(n13350) );
  oai222d1 U1931 ( .A1(n7467), .A2(1'b1), .B1(n12282), .B2(n540), .C1(n7348), 
        .C2(n855), .ZN(n13349) );
  oai222d1 U1930 ( .A1(n7465), .A2(1'b1), .B1(n12281), .B2(n541), .C1(n7342), 
        .C2(n855), .ZN(n13348) );
  oai222d1 U1927 ( .A1(1'b1), .A2(n7445), .B1(n12278), .B2(n541), .C1(n7312), 
        .C2(n855), .ZN(n13345) );
  oai222d1 U1893 ( .A1(1'b1), .A2(n7312), .B1(n12246), .B2(n545), .C1(n876), 
        .C2(n7445), .ZN(n13313) );
  oai222d1 U1955 ( .A1(n7448), .A2(1'b1), .B1(n12306), .B2(n538), .C1(n7318), 
        .C2(n858), .ZN(n13373) );
  oai222d1 U1954 ( .A1(n7438), .A2(1'b1), .B1(n12305), .B2(n538), .C1(n7297), 
        .C2(n858), .ZN(n13372) );
  oai222d1 U1953 ( .A1(n7432), .A2(1'b1), .B1(n12304), .B2(n538), .C1(n7293), 
        .C2(n858), .ZN(n13371) );
  oai222d1 U1952 ( .A1(n7425), .A2(1'b1), .B1(n12303), .B2(n538), .C1(n7288), 
        .C2(n857), .ZN(n13370) );
  oai222d1 U1956 ( .A1(n7514), .A2(1'b1), .B1(n12307), .B2(n538), .C1(n7377), 
        .C2(n858), .ZN(n13374) );
  oai222d1 U1950 ( .A1(n7415), .A2(1'b1), .B1(n12301), .B2(n538), .C1(n7271), 
        .C2(n857), .ZN(n13368) );
  oai222d1 U1949 ( .A1(n7414), .A2(1'b1), .B1(n12300), .B2(n538), .C1(n7265), 
        .C2(n857), .ZN(n13367) );
  oai222d1 U1948 ( .A1(n7412), .A2(1'b1), .B1(n12299), .B2(n539), .C1(n7261), 
        .C2(n857), .ZN(n13366) );
  oai222d1 U1929 ( .A1(n7451), .A2(1'b1), .B1(n12280), .B2(n541), .C1(n7325), 
        .C2(n855), .ZN(n13347) );
  oai222d1 U1928 ( .A1(n7449), .A2(1'b1), .B1(n12279), .B2(n541), .C1(n7322), 
        .C2(n855), .ZN(n13346) );
  oai222d1 U1933 ( .A1(n7476), .A2(1'b1), .B1(n12284), .B2(n540), .C1(n7361), 
        .C2(n855), .ZN(n13351) );
  oai222d1 U1926 ( .A1(n7441), .A2(1'b1), .B1(n12277), .B2(n541), .C1(n7307), 
        .C2(n855), .ZN(n13344) );
  oai222d1 U1892 ( .A1(n7307), .A2(1'b1), .B1(n12245), .B2(n545), .C1(n7441), 
        .C2(n873), .ZN(n13312) );
  oai222d1 U1923 ( .A1(n7408), .A2(1'b1), .B1(n12276), .B2(n542), .C1(n879), 
        .C2(n7558), .ZN(n13343) );
  oai222d1 U1922 ( .A1(n7377), .A2(1'b1), .B1(n12275), .B2(n542), .C1(n879), 
        .C2(n7514), .ZN(n13342) );
  oai222d1 U1921 ( .A1(n7318), .A2(1'b1), .B1(n12274), .B2(n542), .C1(n879), 
        .C2(n7448), .ZN(n13341) );
  oai222d1 U1920 ( .A1(n7297), .A2(1'b1), .B1(n12273), .B2(n542), .C1(n879), 
        .C2(n7438), .ZN(n13340) );
  oai222d1 U2213 ( .A1(n7355), .A2(n788), .B1(n12539), .B2(n777), .C1(n7470), 
        .C2(1'b1), .ZN(n13606) );
  oai222d1 U2214 ( .A1(n7361), .A2(n788), .B1(n12540), .B2(n777), .C1(n7476), 
        .C2(1'b1), .ZN(n13607) );
  oai222d1 U2215 ( .A1(n7363), .A2(n788), .B1(n12541), .B2(n777), .C1(n7482), 
        .C2(1'b1), .ZN(n13608) );
  oai222d1 U2216 ( .A1(n7365), .A2(n788), .B1(n12542), .B2(n777), .C1(n7497), 
        .C2(1'b1), .ZN(n13609) );
  oai222d1 U2217 ( .A1(n7371), .A2(n787), .B1(n12543), .B2(n777), .C1(n7503), 
        .C2(1'b1), .ZN(n13610) );
  oai222d1 U2218 ( .A1(n7372), .A2(n787), .B1(n12544), .B2(n777), .C1(n7510), 
        .C2(1'b1), .ZN(n13611) );
  oai222d1 U2219 ( .A1(n7379), .A2(n787), .B1(n12545), .B2(n777), .C1(n7519), 
        .C2(1'b1), .ZN(n13612) );
  oai222d1 U2220 ( .A1(n7380), .A2(n787), .B1(n12546), .B2(n777), .C1(n7520), 
        .C2(1'b1), .ZN(n13613) );
  oai222d1 U2221 ( .A1(n7387), .A2(n787), .B1(n12547), .B2(n776), .C1(n7524), 
        .C2(1'b1), .ZN(n13614) );
  oai222d1 U2222 ( .A1(n7390), .A2(n787), .B1(n12548), .B2(n776), .C1(n7525), 
        .C2(1'b1), .ZN(n13615) );
  oai222d1 U2223 ( .A1(n7397), .A2(n787), .B1(n12549), .B2(n776), .C1(n7531), 
        .C2(1'b1), .ZN(n13616) );
  oai222d1 U2224 ( .A1(n7398), .A2(n787), .B1(n12550), .B2(n776), .C1(n7538), 
        .C2(1'b1), .ZN(n13617) );
  oai222d1 U2225 ( .A1(n7399), .A2(n787), .B1(n12551), .B2(n776), .C1(n7542), 
        .C2(1'b1), .ZN(n13618) );
  oai222d1 U2226 ( .A1(n7402), .A2(n786), .B1(n12552), .B2(n776), .C1(n7549), 
        .C2(1'b1), .ZN(n13619) );
  oai222d1 U2227 ( .A1(n7403), .A2(n786), .B1(n12553), .B2(n776), .C1(n7552), 
        .C2(1'b1), .ZN(n13620) );
  oai222d1 U2228 ( .A1(n7405), .A2(n786), .B1(n12554), .B2(n776), .C1(n7553), 
        .C2(1'b1), .ZN(n13621) );
  oai222d1 U2229 ( .A1(n7261), .A2(n786), .B1(n12555), .B2(n776), .C1(n7412), 
        .C2(1'b1), .ZN(n13622) );
  oai222d1 U2230 ( .A1(n7265), .A2(n786), .B1(n12556), .B2(n775), .C1(n7414), 
        .C2(1'b1), .ZN(n13623) );
  oai222d1 U1919 ( .A1(n7293), .A2(1'b1), .B1(n12272), .B2(n542), .C1(n879), 
        .C2(n7432), .ZN(n13339) );
  oai222d1 U1918 ( .A1(n7288), .A2(1'b1), .B1(n12271), .B2(n542), .C1(n879), 
        .C2(n7425), .ZN(n13338) );
  oai222d1 U1917 ( .A1(n7278), .A2(1'b1), .B1(n12270), .B2(n542), .C1(n879), 
        .C2(n7424), .ZN(n13337) );
  oai222d1 U1916 ( .A1(n7271), .A2(1'b1), .B1(n12269), .B2(n542), .C1(n879), 
        .C2(n7415), .ZN(n13336) );
  oai222d1 U1915 ( .A1(n7265), .A2(1'b1), .B1(n12268), .B2(n542), .C1(n879), 
        .C2(n7414), .ZN(n13335) );
  oai222d1 U1914 ( .A1(n7261), .A2(1'b1), .B1(n12267), .B2(n543), .C1(n878), 
        .C2(n7412), .ZN(n13334) );
  oai222d1 U1913 ( .A1(n7405), .A2(1'b1), .B1(n12266), .B2(n543), .C1(n878), 
        .C2(n7553), .ZN(n13333) );
  oai222d1 U1912 ( .A1(n7403), .A2(1'b1), .B1(n12265), .B2(n543), .C1(n878), 
        .C2(n7552), .ZN(n13332) );
  oai222d1 U1911 ( .A1(n7402), .A2(1'b1), .B1(n12264), .B2(n543), .C1(n878), 
        .C2(n7549), .ZN(n13331) );
  oai222d1 U1910 ( .A1(n7399), .A2(1'b1), .B1(n12263), .B2(n543), .C1(n878), 
        .C2(n7542), .ZN(n13330) );
  oai222d1 U1909 ( .A1(n7398), .A2(1'b1), .B1(n12262), .B2(n543), .C1(n878), 
        .C2(n7538), .ZN(n13329) );
  oai222d1 U1908 ( .A1(n7397), .A2(1'b1), .B1(n12261), .B2(n543), .C1(n878), 
        .C2(n7531), .ZN(n13328) );
  oai222d1 U1907 ( .A1(n7390), .A2(1'b1), .B1(n12260), .B2(n543), .C1(n878), 
        .C2(n7525), .ZN(n13327) );
  oai222d1 U1906 ( .A1(n7387), .A2(1'b1), .B1(n12259), .B2(n543), .C1(n878), 
        .C2(n7524), .ZN(n13326) );
  oai222d1 U1905 ( .A1(n7380), .A2(1'b1), .B1(n12258), .B2(n544), .C1(n877), 
        .C2(n7520), .ZN(n13325) );
  oai222d1 U1904 ( .A1(n7379), .A2(1'b1), .B1(n12257), .B2(n544), .C1(n877), 
        .C2(n7519), .ZN(n13324) );
  oai222d1 U1903 ( .A1(n7372), .A2(1'b1), .B1(n12256), .B2(n544), .C1(n877), 
        .C2(n7510), .ZN(n13323) );
  oai222d1 U1902 ( .A1(n7371), .A2(1'b1), .B1(n12255), .B2(n544), .C1(n877), 
        .C2(n7503), .ZN(n13322) );
  oai222d1 U1901 ( .A1(n7365), .A2(1'b1), .B1(n12254), .B2(n544), .C1(n877), 
        .C2(n7497), .ZN(n13321) );
  oai222d1 U1900 ( .A1(n7363), .A2(1'b1), .B1(n12253), .B2(n544), .C1(n877), 
        .C2(n7482), .ZN(n13320) );
  oai222d1 U1899 ( .A1(n7361), .A2(1'b1), .B1(n12252), .B2(n544), .C1(n877), 
        .C2(n7476), .ZN(n13319) );
  oai222d1 U1898 ( .A1(n7355), .A2(1'b1), .B1(n12251), .B2(n544), .C1(n877), 
        .C2(n7470), .ZN(n13318) );
  oai222d1 U1897 ( .A1(n7348), .A2(1'b1), .B1(n12250), .B2(n544), .C1(n877), 
        .C2(n7467), .ZN(n13317) );
  oai222d1 U1896 ( .A1(n7342), .A2(1'b1), .B1(n12249), .B2(n545), .C1(n876), 
        .C2(n7465), .ZN(n13316) );
  oai222d1 U1895 ( .A1(n7325), .A2(1'b1), .B1(n12248), .B2(n545), .C1(n876), 
        .C2(n7451), .ZN(n13315) );
  oai222d1 U1894 ( .A1(n7322), .A2(1'b1), .B1(n12247), .B2(n545), .C1(n876), 
        .C2(n7449), .ZN(n13314) );
  oai222d1 U1957 ( .A1(n7558), .A2(1'b1), .B1(n12308), .B2(n538), .C1(n7408), 
        .C2(n858), .ZN(n13375) );
  oai222d1 U2231 ( .A1(n7271), .A2(n786), .B1(n12557), .B2(n775), .C1(n7415), 
        .C2(1'b1), .ZN(n13624) );
  oai222d1 U2232 ( .A1(n7278), .A2(n786), .B1(n12558), .B2(n775), .C1(n7424), 
        .C2(1'b1), .ZN(n13625) );
  oai222d1 U2233 ( .A1(n7288), .A2(n786), .B1(n12559), .B2(n775), .C1(n7425), 
        .C2(1'b1), .ZN(n13626) );
  oai222d1 U2234 ( .A1(n7293), .A2(n786), .B1(n12560), .B2(n775), .C1(n7432), 
        .C2(1'b1), .ZN(n13627) );
  oai222d1 U2235 ( .A1(n7297), .A2(n785), .B1(n12561), .B2(n775), .C1(n7438), 
        .C2(1'b1), .ZN(n13628) );
  oai222d1 U2236 ( .A1(n7318), .A2(n785), .B1(n12562), .B2(n775), .C1(n7448), 
        .C2(1'b1), .ZN(n13629) );
  oai222d1 U2237 ( .A1(n7377), .A2(n785), .B1(n12563), .B2(n775), .C1(n7514), 
        .C2(1'b1), .ZN(n13630) );
  oai222d1 U2238 ( .A1(n7408), .A2(n785), .B1(n12564), .B2(n775), .C1(n7558), 
        .C2(1'b1), .ZN(n13631) );
  oai222d1 U2480 ( .A1(n7432), .A2(n809), .B1(n12528), .B2(n799), .C1(n7293), 
        .C2(1'b1), .ZN(n13792) );
  oai222d1 U2380 ( .A1(n7441), .A2(n721), .B1(n12693), .B2(n717), .C1(n7307), 
        .C2(1'b1), .ZN(n13760) );
  oai222d1 U2383 ( .A1(n7445), .A2(n721), .B1(n12694), .B2(n717), .C1(n7312), 
        .C2(1'b1), .ZN(n13761) );
  oai222d1 U2386 ( .A1(n7449), .A2(n721), .B1(n12695), .B2(n717), .C1(n7322), 
        .C2(1'b1), .ZN(n13762) );
  oai222d1 U2389 ( .A1(n7451), .A2(n721), .B1(n12696), .B2(n717), .C1(n7325), 
        .C2(1'b1), .ZN(n13763) );
  oai222d1 U2392 ( .A1(n7465), .A2(n722), .B1(n12697), .B2(n717), .C1(n7342), 
        .C2(1'b1), .ZN(n13764) );
  oai222d1 U2395 ( .A1(n7467), .A2(n722), .B1(n12698), .B2(n716), .C1(n7348), 
        .C2(1'b1), .ZN(n13765) );
  oai222d1 U2398 ( .A1(n7470), .A2(n722), .B1(n12699), .B2(n716), .C1(n7355), 
        .C2(1'b1), .ZN(n13766) );
  oai222d1 U2401 ( .A1(n7476), .A2(n722), .B1(n12700), .B2(n716), .C1(n7361), 
        .C2(1'b1), .ZN(n13767) );
  oai222d1 U2404 ( .A1(n7482), .A2(n722), .B1(n12701), .B2(n716), .C1(n7363), 
        .C2(1'b1), .ZN(n13768) );
  oai222d1 U2407 ( .A1(n7497), .A2(n722), .B1(n12702), .B2(n716), .C1(n7365), 
        .C2(1'b1), .ZN(n13769) );
  oai222d1 U2410 ( .A1(n7503), .A2(n722), .B1(n12703), .B2(n716), .C1(n7371), 
        .C2(1'b1), .ZN(n13770) );
  oai222d1 U2413 ( .A1(n7510), .A2(n722), .B1(n12704), .B2(n716), .C1(n7372), 
        .C2(1'b1), .ZN(n13771) );
  oai222d1 U2416 ( .A1(n7519), .A2(n722), .B1(n12705), .B2(n716), .C1(n7379), 
        .C2(1'b1), .ZN(n13772) );
  oai222d1 U2419 ( .A1(n7520), .A2(n722), .B1(n12706), .B2(n716), .C1(n7380), 
        .C2(1'b1), .ZN(n13773) );
  oai222d1 U2422 ( .A1(n7524), .A2(n723), .B1(n12707), .B2(n715), .C1(n7387), 
        .C2(1'b1), .ZN(n13774) );
  oai222d1 U2425 ( .A1(n7525), .A2(n723), .B1(n12708), .B2(n715), .C1(n7390), 
        .C2(1'b1), .ZN(n13775) );
  oai222d1 U2428 ( .A1(n7531), .A2(n723), .B1(n12709), .B2(n715), .C1(n7397), 
        .C2(1'b1), .ZN(n13776) );
  oai222d1 U2431 ( .A1(n7538), .A2(n723), .B1(n12710), .B2(n715), .C1(n7398), 
        .C2(1'b1), .ZN(n13777) );
  oai222d1 U2434 ( .A1(n7542), .A2(n723), .B1(n12711), .B2(n715), .C1(n7399), 
        .C2(1'b1), .ZN(n13778) );
  oai222d1 U2437 ( .A1(n7549), .A2(n723), .B1(n12712), .B2(n715), .C1(n7402), 
        .C2(1'b1), .ZN(n13779) );
  oai222d1 U2440 ( .A1(n7552), .A2(n723), .B1(n12713), .B2(n715), .C1(n7403), 
        .C2(1'b1), .ZN(n13780) );
  oai222d1 U2443 ( .A1(n7553), .A2(n723), .B1(n12714), .B2(n715), .C1(n7405), 
        .C2(1'b1), .ZN(n13781) );
  oai222d1 U2446 ( .A1(n7412), .A2(n723), .B1(n12715), .B2(n715), .C1(n7261), 
        .C2(1'b1), .ZN(n13782) );
  oai222d1 U2101 ( .A1(n7441), .A2(n827), .B1(n12437), .B2(n521), .C1(n7307), 
        .C2(1'b1), .ZN(n13504) );
  oai222d1 U2102 ( .A1(n7445), .A2(n827), .B1(n12438), .B2(n521), .C1(n7312), 
        .C2(1'b1), .ZN(n13505) );
  oai222d1 U2103 ( .A1(n7449), .A2(n827), .B1(n12439), .B2(n521), .C1(n7322), 
        .C2(1'b1), .ZN(n13506) );
  oai222d1 U2104 ( .A1(n7451), .A2(n827), .B1(n12440), .B2(n521), .C1(n7325), 
        .C2(1'b1), .ZN(n13507) );
  oai222d1 U2105 ( .A1(n7465), .A2(n828), .B1(n12441), .B2(n521), .C1(n7342), 
        .C2(1'b1), .ZN(n13508) );
  oai222d1 U2106 ( .A1(n7467), .A2(n828), .B1(n12442), .B2(n520), .C1(n7348), 
        .C2(1'b1), .ZN(n13509) );
  oai222d1 U2107 ( .A1(n7470), .A2(n828), .B1(n12443), .B2(n520), .C1(n7355), 
        .C2(1'b1), .ZN(n13510) );
  oai222d1 U2108 ( .A1(n7476), .A2(n828), .B1(n12444), .B2(n520), .C1(n7361), 
        .C2(1'b1), .ZN(n13511) );
  oai222d1 U2109 ( .A1(n7482), .A2(n828), .B1(n12445), .B2(n520), .C1(n7363), 
        .C2(1'b1), .ZN(n13512) );
  oai222d1 U2110 ( .A1(n7497), .A2(n828), .B1(n12446), .B2(n520), .C1(n7365), 
        .C2(1'b1), .ZN(n13513) );
  oai222d1 U2111 ( .A1(n7503), .A2(n828), .B1(n12447), .B2(n520), .C1(n7371), 
        .C2(1'b1), .ZN(n13514) );
  oai222d1 U2112 ( .A1(n7510), .A2(n828), .B1(n12448), .B2(n520), .C1(n7372), 
        .C2(1'b1), .ZN(n13515) );
  oai222d1 U2113 ( .A1(n7519), .A2(n828), .B1(n12449), .B2(n520), .C1(n7379), 
        .C2(1'b1), .ZN(n13516) );
  oai222d1 U2114 ( .A1(n7520), .A2(n828), .B1(n12450), .B2(n520), .C1(n7380), 
        .C2(1'b1), .ZN(n13517) );
  oai222d1 U2115 ( .A1(n7524), .A2(n829), .B1(n12451), .B2(n519), .C1(n7387), 
        .C2(1'b1), .ZN(n13518) );
  oai222d1 U2116 ( .A1(n7525), .A2(n829), .B1(n12452), .B2(n519), .C1(n7390), 
        .C2(1'b1), .ZN(n13519) );
  oai222d1 U2117 ( .A1(n7531), .A2(n829), .B1(n12453), .B2(n519), .C1(n7397), 
        .C2(1'b1), .ZN(n13520) );
  oai222d1 U2118 ( .A1(n7538), .A2(n829), .B1(n12454), .B2(n519), .C1(n7398), 
        .C2(1'b1), .ZN(n13521) );
  oai222d1 U2119 ( .A1(n7542), .A2(n829), .B1(n12455), .B2(n519), .C1(n7399), 
        .C2(1'b1), .ZN(n13522) );
  oai222d1 U2120 ( .A1(n7549), .A2(n829), .B1(n12456), .B2(n519), .C1(n7402), 
        .C2(1'b1), .ZN(n13523) );
  oai222d1 U2121 ( .A1(n7552), .A2(n829), .B1(n12457), .B2(n519), .C1(n7403), 
        .C2(1'b1), .ZN(n13524) );
  oai222d1 U2122 ( .A1(n7553), .A2(n829), .B1(n12458), .B2(n519), .C1(n7405), 
        .C2(1'b1), .ZN(n13525) );
  oai222d1 U2123 ( .A1(n7412), .A2(n829), .B1(n12459), .B2(n519), .C1(n7261), 
        .C2(1'b1), .ZN(n13526) );
  oai222d1 U2124 ( .A1(n7414), .A2(n829), .B1(n12460), .B2(n518), .C1(n7265), 
        .C2(1'b1), .ZN(n13527) );
  oai222d1 U2125 ( .A1(n7415), .A2(n830), .B1(n12461), .B2(n518), .C1(n7271), 
        .C2(1'b1), .ZN(n13528) );
  oai222d1 U2126 ( .A1(n7424), .A2(n830), .B1(n12462), .B2(n518), .C1(n7278), 
        .C2(1'b1), .ZN(n13529) );
  oai222d1 U2127 ( .A1(n7425), .A2(n830), .B1(n12463), .B2(n518), .C1(n7288), 
        .C2(1'b1), .ZN(n13530) );
  oai222d1 U2128 ( .A1(n7432), .A2(n830), .B1(n12464), .B2(n518), .C1(n7293), 
        .C2(1'b1), .ZN(n13531) );
  oai222d1 U2129 ( .A1(n7438), .A2(n830), .B1(n12465), .B2(n518), .C1(n7297), 
        .C2(1'b1), .ZN(n13532) );
  oai222d1 U2130 ( .A1(n7448), .A2(n830), .B1(n12466), .B2(n518), .C1(n7318), 
        .C2(1'b1), .ZN(n13533) );
  oai222d1 U2131 ( .A1(n7514), .A2(n830), .B1(n12467), .B2(n518), .C1(n7377), 
        .C2(1'b1), .ZN(n13534) );
  oai222d1 U2132 ( .A1(n7558), .A2(n830), .B1(n12468), .B2(n518), .C1(n7408), 
        .C2(1'b1), .ZN(n13535) );
  oai222d1 U2449 ( .A1(n7414), .A2(n723), .B1(n12716), .B2(n714), .C1(n7265), 
        .C2(1'b1), .ZN(n13783) );
  oai222d1 U2452 ( .A1(n7415), .A2(n724), .B1(n12717), .B2(n714), .C1(n7271), 
        .C2(1'b1), .ZN(n13784) );
  oai222d1 U2455 ( .A1(n7424), .A2(n724), .B1(n12718), .B2(n714), .C1(n7278), 
        .C2(1'b1), .ZN(n13785) );
  oai222d1 U2458 ( .A1(n7425), .A2(n724), .B1(n12719), .B2(n714), .C1(n7288), 
        .C2(1'b1), .ZN(n13786) );
  oai222d1 U2461 ( .A1(n7432), .A2(n724), .B1(n12720), .B2(n714), .C1(n7293), 
        .C2(1'b1), .ZN(n13787) );
  oai222d1 U2462 ( .A1(n7438), .A2(n724), .B1(n12721), .B2(n714), .C1(n7297), 
        .C2(1'b1), .ZN(n13788) );
  oai222d1 U2465 ( .A1(n7448), .A2(n724), .B1(n12722), .B2(n714), .C1(n7318), 
        .C2(1'b1), .ZN(n13789) );
  oai222d1 U2468 ( .A1(n7514), .A2(n724), .B1(n12723), .B2(n714), .C1(n7377), 
        .C2(1'b1), .ZN(n13790) );
  oai222d1 U2471 ( .A1(n7558), .A2(n724), .B1(n12724), .B2(n714), .C1(n7408), 
        .C2(1'b1), .ZN(n13791) );
  oai222d1 U2141 ( .A1(n7441), .A2(1'b1), .B1(n12469), .B2(n815), .C1(n7307), 
        .C2(n803), .ZN(n13537) );
  oai222d1 U2142 ( .A1(n7445), .A2(1'b1), .B1(n12470), .B2(n815), .C1(n7312), 
        .C2(n803), .ZN(n13538) );
  oai222d1 U2143 ( .A1(n7449), .A2(1'b1), .B1(n12471), .B2(n815), .C1(n7322), 
        .C2(n803), .ZN(n13539) );
  oai222d1 U2144 ( .A1(n7451), .A2(1'b1), .B1(n12472), .B2(n815), .C1(n7325), 
        .C2(n803), .ZN(n13540) );
  oai222d1 U2145 ( .A1(n7465), .A2(1'b1), .B1(n12473), .B2(n815), .C1(n7342), 
        .C2(n803), .ZN(n13541) );
  oai222d1 U2146 ( .A1(n7467), .A2(1'b1), .B1(n12474), .B2(n814), .C1(n7348), 
        .C2(n803), .ZN(n13542) );
  oai222d1 U2147 ( .A1(n7470), .A2(1'b1), .B1(n12475), .B2(n814), .C1(n7355), 
        .C2(n803), .ZN(n13543) );
  oai222d1 U2148 ( .A1(n7476), .A2(1'b1), .B1(n12476), .B2(n814), .C1(n7361), 
        .C2(n803), .ZN(n13544) );
  oai222d1 U2149 ( .A1(n7482), .A2(1'b1), .B1(n12477), .B2(n814), .C1(n7363), 
        .C2(n803), .ZN(n13545) );
  oai222d1 U2150 ( .A1(n7497), .A2(1'b1), .B1(n12478), .B2(n814), .C1(n7365), 
        .C2(n804), .ZN(n13546) );
  oai222d1 U2151 ( .A1(n7503), .A2(1'b1), .B1(n12479), .B2(n814), .C1(n7371), 
        .C2(n804), .ZN(n13547) );
  oai222d1 U2152 ( .A1(n7510), .A2(1'b1), .B1(n12480), .B2(n814), .C1(n7372), 
        .C2(n804), .ZN(n13548) );
  oai222d1 U2153 ( .A1(n7519), .A2(1'b1), .B1(n12481), .B2(n814), .C1(n7379), 
        .C2(n804), .ZN(n13549) );
  oai222d1 U2154 ( .A1(n7520), .A2(1'b1), .B1(n12482), .B2(n814), .C1(n7380), 
        .C2(n804), .ZN(n13550) );
  oai222d1 U2155 ( .A1(n7524), .A2(1'b1), .B1(n12483), .B2(n813), .C1(n7387), 
        .C2(n804), .ZN(n13551) );
  oai222d1 U2156 ( .A1(n7525), .A2(1'b1), .B1(n12484), .B2(n813), .C1(n7390), 
        .C2(n804), .ZN(n13552) );
  oai222d1 U2157 ( .A1(n7531), .A2(1'b1), .B1(n12485), .B2(n813), .C1(n7397), 
        .C2(n804), .ZN(n13553) );
  oai222d1 U2158 ( .A1(n7538), .A2(1'b1), .B1(n12486), .B2(n813), .C1(n7398), 
        .C2(n804), .ZN(n13554) );
  oai222d1 U2159 ( .A1(n7542), .A2(1'b1), .B1(n12487), .B2(n813), .C1(n7399), 
        .C2(n805), .ZN(n13555) );
  oai222d1 U2160 ( .A1(n7549), .A2(1'b1), .B1(n12488), .B2(n813), .C1(n7402), 
        .C2(n805), .ZN(n13556) );
  oai222d1 U2161 ( .A1(n7552), .A2(1'b1), .B1(n12489), .B2(n813), .C1(n7403), 
        .C2(n805), .ZN(n13557) );
  oai222d1 U2162 ( .A1(n7553), .A2(1'b1), .B1(n12490), .B2(n813), .C1(n7405), 
        .C2(n805), .ZN(n13558) );
  oai222d1 U2163 ( .A1(n7412), .A2(1'b1), .B1(n12491), .B2(n813), .C1(n7261), 
        .C2(n805), .ZN(n13559) );
  oai222d1 U1861 ( .A1(1'b1), .A2(n7441), .B1(n12213), .B2(n517), .C1(n876), 
        .C2(n7307), .ZN(n13281) );
  oai222d1 U1862 ( .A1(1'b1), .A2(n7449), .B1(n12215), .B2(n517), .C1(n873), 
        .C2(n7322), .ZN(n13282) );
  oai222d1 U1863 ( .A1(1'b1), .A2(n7451), .B1(n12216), .B2(n517), .C1(n873), 
        .C2(n7325), .ZN(n13283) );
  oai222d1 U1864 ( .A1(1'b1), .A2(n7465), .B1(n12217), .B2(n517), .C1(n873), 
        .C2(n7342), .ZN(n13284) );
  oai222d1 U1865 ( .A1(1'b1), .A2(n7467), .B1(n12218), .B2(n517), .C1(n873), 
        .C2(n7348), .ZN(n13285) );
  oai222d1 U1866 ( .A1(1'b1), .A2(n7470), .B1(n12219), .B2(n516), .C1(n873), 
        .C2(n7355), .ZN(n13286) );
  oai222d1 U1867 ( .A1(1'b1), .A2(n7476), .B1(n12220), .B2(n516), .C1(n873), 
        .C2(n7361), .ZN(n13287) );
  oai222d1 U1868 ( .A1(1'b1), .A2(n7482), .B1(n12221), .B2(n516), .C1(n873), 
        .C2(n7363), .ZN(n13288) );
  oai222d1 U1869 ( .A1(1'b1), .A2(n7497), .B1(n12222), .B2(n516), .C1(n873), 
        .C2(n7365), .ZN(n13289) );
  oai222d1 U1870 ( .A1(1'b1), .A2(n7503), .B1(n12223), .B2(n516), .C1(n874), 
        .C2(n7371), .ZN(n13290) );
  oai222d1 U1871 ( .A1(1'b1), .A2(n7510), .B1(n12224), .B2(n516), .C1(n874), 
        .C2(n7372), .ZN(n13291) );
  oai222d1 U1872 ( .A1(1'b1), .A2(n7519), .B1(n12225), .B2(n516), .C1(n874), 
        .C2(n7379), .ZN(n13292) );
  oai222d1 U1873 ( .A1(1'b1), .A2(n7520), .B1(n12226), .B2(n516), .C1(n874), 
        .C2(n7380), .ZN(n13293) );
  oai222d1 U1874 ( .A1(1'b1), .A2(n7524), .B1(n12227), .B2(n516), .C1(n874), 
        .C2(n7387), .ZN(n13294) );
  oai222d1 U1875 ( .A1(1'b1), .A2(n7525), .B1(n12228), .B2(n515), .C1(n874), 
        .C2(n7390), .ZN(n13295) );
  oai222d1 U1876 ( .A1(1'b1), .A2(n7531), .B1(n12229), .B2(n515), .C1(n874), 
        .C2(n7397), .ZN(n13296) );
  oai222d1 U1877 ( .A1(1'b1), .A2(n7538), .B1(n12230), .B2(n515), .C1(n874), 
        .C2(n7398), .ZN(n13297) );
  oai222d1 U1878 ( .A1(1'b1), .A2(n7542), .B1(n12231), .B2(n515), .C1(n874), 
        .C2(n7399), .ZN(n13298) );
  oai222d1 U1879 ( .A1(1'b1), .A2(n7549), .B1(n12232), .B2(n515), .C1(n875), 
        .C2(n7402), .ZN(n13299) );
  oai222d1 U1880 ( .A1(1'b1), .A2(n7552), .B1(n12233), .B2(n515), .C1(n875), 
        .C2(n7403), .ZN(n13300) );
  oai222d1 U1881 ( .A1(1'b1), .A2(n7553), .B1(n12234), .B2(n515), .C1(n875), 
        .C2(n7405), .ZN(n13301) );
  oai222d1 U1882 ( .A1(1'b1), .A2(n7412), .B1(n12235), .B2(n515), .C1(n875), 
        .C2(n7261), .ZN(n13302) );
  oai222d1 U1883 ( .A1(1'b1), .A2(n7414), .B1(n12236), .B2(n515), .C1(n875), 
        .C2(n7265), .ZN(n13303) );
  oai222d1 U1884 ( .A1(1'b1), .A2(n7415), .B1(n12237), .B2(n514), .C1(n875), 
        .C2(n7271), .ZN(n13304) );
  oai222d1 U1885 ( .A1(1'b1), .A2(n7424), .B1(n12238), .B2(n514), .C1(n875), 
        .C2(n7278), .ZN(n13305) );
  oai222d1 U1886 ( .A1(1'b1), .A2(n7425), .B1(n12239), .B2(n514), .C1(n875), 
        .C2(n7288), .ZN(n13306) );
  oai222d1 U1887 ( .A1(1'b1), .A2(n7432), .B1(n12240), .B2(n514), .C1(n875), 
        .C2(n7293), .ZN(n13307) );
  oai222d1 U1888 ( .A1(1'b1), .A2(n7438), .B1(n12241), .B2(n514), .C1(n876), 
        .C2(n7297), .ZN(n13308) );
  oai222d1 U1889 ( .A1(1'b1), .A2(n7448), .B1(n12242), .B2(n514), .C1(n876), 
        .C2(n7318), .ZN(n13309) );
  oai222d1 U1890 ( .A1(1'b1), .A2(n7514), .B1(n12243), .B2(n514), .C1(n876), 
        .C2(n7377), .ZN(n13310) );
  oai222d1 U1891 ( .A1(1'b1), .A2(n7558), .B1(n12244), .B2(n514), .C1(n876), 
        .C2(n7408), .ZN(n13311) );
  oai222d1 U2137 ( .A1(1'b1), .A2(n7445), .B1(n12214), .B2(n514), .C1(n880), 
        .C2(n7312), .ZN(n13536) );
  oai222d1 U2164 ( .A1(n7414), .A2(1'b1), .B1(n12492), .B2(n812), .C1(n7265), 
        .C2(n805), .ZN(n13560) );
  oai222d1 U2165 ( .A1(n7415), .A2(1'b1), .B1(n12493), .B2(n812), .C1(n7271), 
        .C2(n805), .ZN(n13561) );
  oai222d1 U2166 ( .A1(n7424), .A2(1'b1), .B1(n12494), .B2(n812), .C1(n7278), 
        .C2(n805), .ZN(n13562) );
  oai222d1 U2167 ( .A1(n7425), .A2(1'b1), .B1(n12495), .B2(n812), .C1(n7288), 
        .C2(n805), .ZN(n13563) );
  oai222d1 U2168 ( .A1(n7432), .A2(1'b1), .B1(n12496), .B2(n812), .C1(n7293), 
        .C2(n806), .ZN(n13564) );
  oai222d1 U2169 ( .A1(n7438), .A2(1'b1), .B1(n12497), .B2(n812), .C1(n7297), 
        .C2(n806), .ZN(n13565) );
  oai222d1 U2170 ( .A1(n7448), .A2(1'b1), .B1(n12498), .B2(n812), .C1(n7318), 
        .C2(n806), .ZN(n13566) );
  oai222d1 U2171 ( .A1(n7514), .A2(1'b1), .B1(n12499), .B2(n812), .C1(n7377), 
        .C2(n806), .ZN(n13567) );
  oai222d1 U2172 ( .A1(n7558), .A2(1'b1), .B1(n12500), .B2(n812), .C1(n7408), 
        .C2(n806), .ZN(n13568) );
  invbd2 U4 ( .I(n4355), .ZN(N26480) );
  aoi211d1 U5 ( .C1(1'b1), .C2(n954), .A(n1), .B(n3583), .ZN(n3581) );
  invbd2 U6 ( .I(n949), .ZN(n3580) );
  invbd2 U8 ( .I(n3620), .ZN(n12105) );
  nd02d2 U9 ( .A1(reorder_A1[0]), .A2(n3623), .ZN(n3620) );
  nr02d2 U10 ( .A1(N3855), .A2(n2788), .ZN(n4362) );
  nd02d2 U11 ( .A1(n2781), .A2(n495), .ZN(n4350) );
  nd02d2 U12 ( .A1(n4345), .A2(n495), .ZN(n4349) );
  nd02d2 U13 ( .A1(n4337), .A2(n495), .ZN(n4340) );
  nd02d2 U14 ( .A1(n4345), .A2(n495), .ZN(n4344) );
  nd02d2 U17 ( .A1(n4329), .A2(n495), .ZN(n4332) );
  nd02d2 U20 ( .A1(n4337), .A2(n495), .ZN(n4336) );
  nr02d1 U21 ( .A1(n14), .A2(n7882), .ZN(n7889) );
  nr02d1 U22 ( .A1(n20), .A2(n9376), .ZN(n11737) );
  nr02d1 U23 ( .A1(n26), .A2(n5321), .ZN(n10407) );
  an03d1 U24 ( .A1(n3647), .A2(n2770), .A3(n3651), .Z(n1) );
  nr02d1 U25 ( .A1(n3667), .A2(n3656), .ZN(n2) );
  an02d1 U26 ( .A1(n417), .A2(n485), .Z(n3) );
  or02d1 U27 ( .A1(n1853), .A2(n1370), .Z(n4) );
  aor211d1 U28 ( .C1(n1014), .C2(n968), .A(n2624), .B(n12), .Z(n5) );
  nr02d1 U29 ( .A1(\sub_183/carry[8] ), .A2(n1340), .ZN(n6) );
  buffd1 U30 ( .I(n1218), .Z(n1217) );
  buffd1 U31 ( .I(n1320), .Z(n1318) );
  buffd1 U32 ( .I(n1129), .Z(n1128) );
  buffd1 U33 ( .I(n1321), .Z(n1317) );
  buffd1 U34 ( .I(n1321), .Z(n1315) );
  buffd1 U35 ( .I(n1268), .Z(n1260) );
  buffd1 U36 ( .I(n1321), .Z(n1316) );
  buffd1 U37 ( .I(n1322), .Z(n1313) );
  buffd1 U38 ( .I(n1268), .Z(n1261) );
  buffd1 U39 ( .I(n1130), .Z(n1125) );
  buffd1 U40 ( .I(n1174), .Z(n1164) );
  buffd1 U41 ( .I(n1268), .Z(n1259) );
  buffd1 U42 ( .I(n1267), .Z(n1263) );
  buffd1 U43 ( .I(n1219), .Z(n1215) );
  buffd1 U44 ( .I(n1220), .Z(n1212) );
  buffd1 U45 ( .I(n1219), .Z(n1214) );
  buffd1 U46 ( .I(n1322), .Z(n1312) );
  buffd1 U47 ( .I(n1220), .Z(n1211) );
  buffd1 U48 ( .I(n1220), .Z(n1210) );
  buffd1 U49 ( .I(n1267), .Z(n1264) );
  buffd1 U50 ( .I(n1174), .Z(n1165) );
  buffd1 U51 ( .I(n1173), .Z(n1168) );
  buffd1 U52 ( .I(n1173), .Z(n1169) );
  buffd1 U53 ( .I(n1129), .Z(n1126) );
  buffd1 U54 ( .I(n1130), .Z(n1123) );
  buffd1 U55 ( .I(n1173), .Z(n1167) );
  buffd1 U56 ( .I(n1129), .Z(n1127) );
  buffd1 U57 ( .I(n1174), .Z(n1166) );
  buffd1 U58 ( .I(n1130), .Z(n1124) );
  buffd1 U59 ( .I(n1218), .Z(n1216) );
  buffd1 U60 ( .I(n1172), .Z(n1170) );
  buffd1 U61 ( .I(n1266), .Z(n1265) );
  buffd1 U62 ( .I(n1131), .Z(n1122) );
  buffd1 U63 ( .I(n1323), .Z(n1310) );
  buffd1 U64 ( .I(n1323), .Z(n1311) );
  buffd1 U65 ( .I(n1371), .Z(n1353) );
  buffd1 U66 ( .I(n1370), .Z(n1356) );
  buffd1 U67 ( .I(n1370), .Z(n1354) );
  buffd1 U68 ( .I(n1371), .Z(n1352) );
  buffd1 U69 ( .I(n1370), .Z(n1355) );
  buffd1 U70 ( .I(n1371), .Z(n1351) );
  buffd1 U71 ( .I(n1267), .Z(n1262) );
  buffd1 U72 ( .I(n1322), .Z(n1314) );
  buffd1 U73 ( .I(n1219), .Z(n1213) );
  buffd1 U74 ( .I(n1131), .Z(n1121) );
  buffd1 U75 ( .I(n1036), .Z(n1031) );
  buffd1 U76 ( .I(n1036), .Z(n1032) );
  buffd1 U77 ( .I(n1036), .Z(n1030) );
  buffd1 U78 ( .I(n1036), .Z(n1029) );
  buffd1 U79 ( .I(n1036), .Z(n1033) );
  buffd1 U80 ( .I(n1269), .Z(n1258) );
  inv0d0 U81 ( .I(N3972), .ZN(n512) );
  inv0d0 U82 ( .I(N3974), .ZN(n501) );
  inv0d0 U83 ( .I(N3973), .ZN(n499) );
  inv0d0 U84 ( .I(N3179), .ZN(n505) );
  inv0d0 U85 ( .I(N3976), .ZN(n503) );
  inv0d0 U86 ( .I(N3180), .ZN(n507) );
  inv0d0 U87 ( .I(N3975), .ZN(n956) );
  inv0d0 U88 ( .I(N3855), .ZN(n511) );
  inv0d0 U89 ( .I(num_images[1]), .ZN(n1036) );
  inv0d0 U90 ( .I(n1222), .ZN(n1221) );
  inv0d0 U91 ( .I(n1271), .ZN(n1270) );
  inv0d0 U92 ( .I(n958), .ZN(n957) );
  inv0d0 U93 ( .I(n1088), .ZN(n1087) );
  inv0d0 U94 ( .I(n1133), .ZN(n1132) );
  inv0d0 U95 ( .I(n1176), .ZN(n1175) );
  inv0d0 U96 ( .I(n5565), .ZN(n3028) );
  nd02d1 U97 ( .A1(n3034), .A2(n3029), .ZN(n5565) );
  inv0d0 U98 ( .I(n8725), .ZN(n3095) );
  inv0d0 U99 ( .I(n7534), .ZN(n4188) );
  inv0d0 U100 ( .I(n10129), .ZN(n3171) );
  inv0d0 U101 ( .I(n7783), .ZN(n3429) );
  inv0d0 U102 ( .I(n4403), .ZN(n4028) );
  inv0d0 U103 ( .I(n485), .ZN(n486) );
  buffd1 U104 ( .I(n466), .Z(n461) );
  buffd1 U105 ( .I(n465), .Z(n458) );
  buffd1 U106 ( .I(n467), .Z(n462) );
  buffd1 U107 ( .I(n466), .Z(n459) );
  buffd1 U108 ( .I(n475), .Z(n471) );
  buffd1 U109 ( .I(n476), .Z(n468) );
  buffd1 U110 ( .I(n467), .Z(n463) );
  buffd1 U111 ( .I(n476), .Z(n472) );
  buffd1 U112 ( .I(n475), .Z(n469) );
  buffd1 U113 ( .I(n466), .Z(n460) );
  buffd1 U114 ( .I(n467), .Z(n464) );
  buffd1 U115 ( .I(n476), .Z(n473) );
  buffd1 U116 ( .I(n475), .Z(n470) );
  buffd1 U117 ( .I(n476), .Z(n474) );
  buffd1 U118 ( .I(n481), .Z(n479) );
  buffd1 U119 ( .I(n480), .Z(n477) );
  buffd1 U120 ( .I(n480), .Z(n478) );
  inv0d0 U121 ( .I(n4757), .ZN(n3090) );
  inv0d0 U122 ( .I(n5396), .ZN(n3465) );
  nd02d1 U123 ( .A1(n4191), .A2(n4189), .ZN(n7534) );
  nd02d1 U124 ( .A1(n3372), .A2(n3413), .ZN(n4547) );
  nd02d1 U125 ( .A1(n3463), .A2(n3431), .ZN(n7783) );
  inv0d0 U126 ( .I(n4929), .ZN(n2828) );
  nd02d1 U127 ( .A1(n6854), .A2(n4053), .ZN(n4403) );
  nd02d1 U128 ( .A1(n3097), .A2(n3108), .ZN(n8725) );
  inv0d0 U129 ( .I(n6092), .ZN(n3801) );
  inv0d0 U130 ( .I(n4803), .ZN(n2955) );
  inv0d0 U131 ( .I(n1378), .ZN(n1380) );
  inv0d0 U132 ( .I(n5076), .ZN(n4053) );
  inv0d0 U133 ( .I(n4713), .ZN(n3041) );
  inv0d0 U134 ( .I(n4744), .ZN(n3073) );
  nd02d1 U135 ( .A1(n3173), .A2(n3174), .ZN(n10129) );
  inv0d0 U136 ( .I(n4704), .ZN(n3029) );
  inv0d0 U137 ( .I(n10279), .ZN(n2842) );
  inv0d0 U138 ( .I(n2576), .ZN(n2578) );
  inv0d0 U139 ( .I(n8057), .ZN(n3223) );
  inv0d0 U140 ( .I(n2555), .ZN(n2556) );
  inv0d0 U141 ( .I(n4876), .ZN(n2869) );
  inv0d0 U142 ( .I(n5597), .ZN(n3072) );
  inv0d0 U143 ( .I(n12068), .ZN(n4178) );
  inv0d0 U144 ( .I(n6978), .ZN(n3751) );
  inv0d0 U145 ( .I(n2326), .ZN(n2328) );
  inv0d0 U146 ( .I(n7344), .ZN(n2850) );
  inv0d0 U147 ( .I(n8774), .ZN(n2976) );
  inv0d0 U148 ( .I(n6434), .ZN(n3034) );
  inv0d0 U149 ( .I(n8235), .ZN(n4191) );
  inv0d0 U150 ( .I(n5654), .ZN(n2989) );
  inv0d0 U151 ( .I(n4390), .ZN(n3822) );
  inv0d0 U152 ( .I(n10198), .ZN(n3081) );
  inv0d0 U153 ( .I(n7970), .ZN(n3015) );
  inv0d0 U154 ( .I(n9445), .ZN(n3218) );
  inv0d0 U155 ( .I(n9447), .ZN(n3216) );
  inv0d0 U156 ( .I(n8056), .ZN(n3215) );
  inv0d0 U157 ( .I(n1524), .ZN(n1525) );
  inv0d0 U158 ( .I(n2111), .ZN(n2112) );
  inv0d0 U159 ( .I(n2119), .ZN(n2120) );
  inv0d0 U160 ( .I(n1491), .ZN(n1492) );
  inv0d0 U161 ( .I(n1499), .ZN(n1500) );
  inv0d0 U162 ( .I(n4655), .ZN(n3174) );
  inv0d0 U163 ( .I(n8295), .ZN(n4081) );
  inv0d0 U164 ( .I(n2126), .ZN(n2127) );
  inv0d0 U165 ( .I(n9490), .ZN(n3100) );
  inv0d0 U166 ( .I(n5393), .ZN(n3463) );
  inv0d0 U167 ( .I(n4856), .ZN(n2826) );
  inv0d0 U168 ( .I(n5028), .ZN(n4072) );
  inv0d0 U169 ( .I(n11602), .ZN(n3668) );
  inv0d0 U170 ( .I(n10874), .ZN(n3374) );
  inv0d0 U171 ( .I(n5347), .ZN(n3574) );
  inv0d0 U172 ( .I(n7644), .ZN(n4032) );
  inv0d0 U173 ( .I(n5169), .ZN(n3970) );
  inv0d0 U174 ( .I(n5066), .ZN(n4017) );
  inv0d0 U175 ( .I(n4971), .ZN(n3164) );
  inv0d0 U176 ( .I(n5661), .ZN(n2959) );
  buffd1 U177 ( .I(n10), .Z(n485) );
  inv0d0 U178 ( .I(n483), .ZN(n489) );
  inv0d0 U179 ( .I(n482), .ZN(n490) );
  inv0d0 U180 ( .I(n484), .ZN(n487) );
  buffd1 U181 ( .I(n10), .Z(n484) );
  inv0d0 U182 ( .I(n483), .ZN(n491) );
  buffd1 U183 ( .I(n10), .Z(n483) );
  inv0d0 U184 ( .I(n484), .ZN(n488) );
  inv0d0 U185 ( .I(n482), .ZN(n492) );
  buffd1 U186 ( .I(n10), .Z(n482) );
  buffd1 U187 ( .I(n428), .Z(n423) );
  buffd1 U188 ( .I(n427), .Z(n420) );
  buffd1 U189 ( .I(n395), .Z(n466) );
  buffd1 U190 ( .I(n395), .Z(n465) );
  buffd1 U191 ( .I(n429), .Z(n424) );
  buffd1 U192 ( .I(n428), .Z(n421) );
  buffd1 U193 ( .I(n395), .Z(n467) );
  buffd1 U194 ( .I(n437), .Z(n433) );
  buffd1 U195 ( .I(n447), .Z(n442) );
  buffd1 U196 ( .I(n438), .Z(n430) );
  buffd1 U197 ( .I(n446), .Z(n439) );
  buffd1 U198 ( .I(n396), .Z(n475) );
  buffd1 U199 ( .I(n429), .Z(n425) );
  buffd1 U200 ( .I(n438), .Z(n434) );
  buffd1 U201 ( .I(n437), .Z(n431) );
  buffd1 U202 ( .I(n448), .Z(n443) );
  buffd1 U203 ( .I(n447), .Z(n440) );
  buffd1 U204 ( .I(n396), .Z(n476) );
  buffd1 U205 ( .I(n428), .Z(n422) );
  buffd1 U206 ( .I(n456), .Z(n452) );
  buffd1 U207 ( .I(n429), .Z(n426) );
  buffd1 U208 ( .I(n457), .Z(n449) );
  buffd1 U209 ( .I(n438), .Z(n435) );
  buffd1 U210 ( .I(n448), .Z(n444) );
  buffd1 U211 ( .I(n457), .Z(n453) );
  buffd1 U212 ( .I(n456), .Z(n450) );
  buffd1 U213 ( .I(n437), .Z(n432) );
  buffd1 U214 ( .I(n438), .Z(n436) );
  buffd1 U215 ( .I(n447), .Z(n441) );
  buffd1 U216 ( .I(n448), .Z(n445) );
  buffd1 U217 ( .I(n397), .Z(n481) );
  buffd1 U218 ( .I(n457), .Z(n454) );
  buffd1 U219 ( .I(n397), .Z(n480) );
  buffd1 U220 ( .I(n456), .Z(n451) );
  buffd1 U221 ( .I(n457), .Z(n455) );
  inv0d0 U222 ( .I(n3617), .ZN(n2754) );
  buffd1 U223 ( .I(n870), .Z(n873) );
  buffd1 U224 ( .I(n871), .Z(n878) );
  buffd1 U225 ( .I(n871), .Z(n877) );
  buffd1 U226 ( .I(n870), .Z(n875) );
  buffd1 U227 ( .I(n870), .Z(n874) );
  buffd1 U228 ( .I(n871), .Z(n876) );
  buffd1 U229 ( .I(n872), .Z(n879) );
  buffd1 U230 ( .I(n872), .Z(n880) );
  nd02d1 U231 ( .A1(N12226), .A2(n3467), .ZN(n5396) );
  nd02d1 U232 ( .A1(n2829), .A2(n2849), .ZN(n4929) );
  nd03d1 U233 ( .A1(n3850), .A2(n3851), .A3(n3955), .ZN(n4400) );
  inv0d0 U234 ( .I(n2149), .ZN(n2151) );
  nr02d1 U235 ( .A1(n6588), .A2(n8057), .ZN(n9447) );
  nd02d1 U236 ( .A1(n3045), .A2(n3043), .ZN(n4713) );
  nd02d1 U237 ( .A1(n3231), .A2(n3224), .ZN(n8057) );
  nd02d1 U238 ( .A1(n2956), .A2(n3004), .ZN(n4803) );
  nr02d1 U239 ( .A1(n4872), .A2(n2871), .ZN(n4878) );
  nr02d1 U240 ( .A1(n3314), .A2(n3282), .ZN(n5486) );
  nd02d1 U241 ( .A1(n2979), .A2(n2980), .ZN(n8774) );
  inv0d0 U242 ( .I(n1674), .ZN(n1677) );
  inv0d0 U243 ( .I(n1826), .ZN(n1829) );
  nd02d1 U244 ( .A1(N9876), .A2(n4054), .ZN(n5076) );
  nd02d1 U245 ( .A1(n3121), .A2(n3073), .ZN(n5597) );
  nd02d1 U246 ( .A1(n3030), .A2(n3227), .ZN(n4704) );
  nd02d1 U247 ( .A1(n3823), .A2(n3832), .ZN(n4390) );
  nd02d1 U248 ( .A1(n3759), .A2(n3757), .ZN(n6978) );
  nd02d1 U249 ( .A1(n3275), .A2(n3330), .ZN(n5475) );
  nd02d1 U250 ( .A1(n4018), .A2(n10603), .ZN(n5066) );
  nd02d1 U251 ( .A1(n4063), .A2(n4116), .ZN(n5882) );
  nd02d1 U252 ( .A1(n3016), .A2(n5619), .ZN(n7970) );
  nr02d1 U253 ( .A1(n10613), .A2(n5095), .ZN(n6854) );
  nd02d1 U254 ( .A1(n4810), .A2(n2990), .ZN(n5654) );
  nr02d1 U255 ( .A1(n4407), .A2(n6978), .ZN(n7718) );
  nd02d1 U256 ( .A1(n4104), .A2(n4108), .ZN(n5026) );
  nd02d1 U257 ( .A1(n3971), .A2(n5093), .ZN(n5169) );
  nd02d1 U258 ( .A1(n3089), .A2(n4764), .ZN(n5616) );
  nd02d1 U259 ( .A1(n3075), .A2(n3074), .ZN(n4744) );
  nd02d1 U260 ( .A1(n3199), .A2(n3241), .ZN(n4671) );
  nd02d1 U261 ( .A1(n3248), .A2(n3250), .ZN(n4638) );
  nr02d1 U262 ( .A1(n7534), .A2(n5810), .ZN(n7530) );
  nd12d1 U263 ( .A1(n7), .A2(n2849), .ZN(n10279) );
  nd04d1 U264 ( .A1(n1343), .A2(n1299), .A3(n1246), .A4(n1200), .ZN(n7) );
  nd02d1 U265 ( .A1(n4160), .A2(n4175), .ZN(n5853) );
  nd02d1 U266 ( .A1(n3920), .A2(n6883), .ZN(n6880) );
  inv0d0 U267 ( .I(n4810), .ZN(n2999) );
  nd02d1 U268 ( .A1(n5678), .A2(n2828), .ZN(n4856) );
  nd02d1 U269 ( .A1(n2870), .A2(n2871), .ZN(n4876) );
  inv0d0 U270 ( .I(n11071), .ZN(n3097) );
  nd02d1 U271 ( .A1(n8807), .A2(n2878), .ZN(n4884) );
  nd02d1 U272 ( .A1(n3094), .A2(n9599), .ZN(n4757) );
  nd03d1 U273 ( .A1(n3299), .A2(n3294), .A3(n3165), .ZN(n4971) );
  nd02d1 U274 ( .A1(n3464), .A2(n3465), .ZN(n5393) );
  nd02d1 U275 ( .A1(n4196), .A2(n4195), .ZN(n8235) );
  nd02d1 U276 ( .A1(n2968), .A2(n2962), .ZN(n5661) );
  nd02d1 U277 ( .A1(N11316), .A2(n3802), .ZN(n6092) );
  nd02d1 U278 ( .A1(N9966), .A2(n4049), .ZN(n5095) );
  nd02d1 U279 ( .A1(n2944), .A2(n4798), .ZN(n5641) );
  nd02d1 U280 ( .A1(n3179), .A2(n3175), .ZN(n4655) );
  nd02d1 U281 ( .A1(n3037), .A2(n3035), .ZN(n6434) );
  nd02d1 U282 ( .A1(n9554), .A2(n2913), .ZN(n7344) );
  nd02d1 U283 ( .A1(n3041), .A2(n3037), .ZN(n8675) );
  nd02d1 U284 ( .A1(n5619), .A2(n4764), .ZN(n9490) );
  nd02d1 U285 ( .A1(n4073), .A2(n4110), .ZN(n5028) );
  inv0d0 U286 ( .I(n6465), .ZN(n3065) );
  nd02d1 U287 ( .A1(n3575), .A2(n3788), .ZN(n5347) );
  inv0d0 U288 ( .I(n8307), .ZN(n3998) );
  inv0d0 U289 ( .I(n8722), .ZN(n3108) );
  inv0d0 U290 ( .I(n8534), .ZN(n3456) );
  inv0d0 U291 ( .I(n6316), .ZN(n3282) );
  or03d0 U292 ( .A1(n1307), .A2(n1233), .A3(n1183), .Z(n8) );
  inv0d0 U293 ( .I(N8008), .ZN(n7574) );
  inv0d0 U294 ( .I(n5287), .ZN(n3742) );
  inv0d0 U295 ( .I(n4721), .ZN(n3047) );
  nd02d1 U296 ( .A1(n6316), .A2(n3313), .ZN(n4607) );
  nd12d1 U297 ( .A1(n9), .A2(n4179), .ZN(n12068) );
  aoi211d1 U298 ( .C1(n1239), .C2(n2503), .A(n1339), .B(n1280), .ZN(n9) );
  nd02d1 U299 ( .A1(n9447), .A2(n3211), .ZN(n7247) );
  nd03d1 U300 ( .A1(n9957), .A2(n3798), .A3(n3769), .ZN(n8449) );
  nd02d1 U301 ( .A1(n3326), .A2(n3323), .ZN(n5478) );
  inv0d0 U302 ( .I(n9202), .ZN(n3757) );
  nd02d1 U303 ( .A1(n3909), .A2(n3911), .ZN(n4418) );
  inv0d0 U304 ( .I(n7331), .ZN(n2979) );
  inv0d0 U305 ( .I(n8787), .ZN(n2845) );
  nd02d1 U306 ( .A1(n3401), .A2(n3375), .ZN(n10874) );
  inv0d0 U307 ( .I(n6691), .ZN(n4238) );
  nd02d1 U308 ( .A1(n4038), .A2(n4033), .ZN(n7644) );
  nd02d1 U309 ( .A1(n2978), .A2(n4933), .ZN(n4846) );
  nd02d1 U310 ( .A1(n3117), .A2(n3084), .ZN(n10198) );
  inv0d0 U311 ( .I(n4545), .ZN(n3413) );
  nd02d1 U312 ( .A1(n3316), .A2(n3319), .ZN(n9388) );
  nd02d1 U313 ( .A1(n11003), .A2(n3223), .ZN(n8056) );
  inv0d0 U314 ( .I(n4696), .ZN(n3027) );
  nd02d1 U315 ( .A1(n4082), .A2(n4104), .ZN(n8295) );
  nd02d1 U316 ( .A1(n3738), .A2(n3751), .ZN(n4401) );
  nd02d1 U317 ( .A1(n3573), .A2(n3575), .ZN(n8077) );
  nd02d1 U318 ( .A1(n2888), .A2(n2894), .ZN(n4908) );
  nd02d1 U319 ( .A1(n2893), .A2(n2888), .ZN(n4906) );
  nd02d1 U320 ( .A1(n3672), .A2(n4692), .ZN(n11602) );
  nd02d1 U321 ( .A1(n3227), .A2(n3219), .ZN(n9445) );
  inv0d0 U322 ( .I(n9562), .ZN(n2876) );
  nd02d1 U323 ( .A1(n3957), .A2(n3819), .ZN(n6009) );
  nd02d1 U324 ( .A1(n10942), .A2(n5505), .ZN(n9401) );
  nd02d1 U325 ( .A1(n4279), .A2(n4281), .ZN(n8179) );
  nd02d1 U326 ( .A1(n7287), .A2(n9599), .ZN(n6474) );
  inv0d0 U327 ( .I(n5402), .ZN(n3431) );
  inv0d0 U328 ( .I(n6203), .ZN(n3367) );
  inv0d0 U329 ( .I(n11623), .ZN(n3788) );
  inv0d0 U330 ( .I(n10674), .ZN(n3836) );
  inv0d0 U331 ( .I(n4739), .ZN(n3064) );
  inv0d0 U332 ( .I(n6063), .ZN(n3730) );
  inv0d0 U333 ( .I(N8107), .ZN(n7588) );
  inv0d0 U334 ( .I(n8171), .ZN(n4376) );
  inv0d0 U335 ( .I(n4586), .ZN(n3326) );
  inv0d0 U336 ( .I(n6616), .ZN(n3537) );
  inv0d0 U337 ( .I(n4715), .ZN(n3046) );
  inv0d0 U338 ( .I(n6528), .ZN(n2961) );
  inv0d0 U339 ( .I(n2542), .ZN(n2546) );
  inv0d0 U340 ( .I(n7614), .ZN(n4016) );
  inv0d0 U341 ( .I(n5445), .ZN(n3405) );
  inv0d0 U342 ( .I(n7747), .ZN(n3521) );
  inv0d0 U343 ( .I(n8622), .ZN(n3175) );
  inv0d0 U344 ( .I(n9185), .ZN(n3862) );
  inv0d0 U345 ( .I(n7139), .ZN(n3387) );
  inv0d0 U346 ( .I(n11803), .ZN(n3204) );
  inv0d0 U347 ( .I(n4779), .ZN(n2926) );
  inv0d0 U348 ( .I(n5619), .ZN(n3099) );
  inv0d0 U349 ( .I(n5805), .ZN(n4189) );
  inv0d0 U350 ( .I(n7059), .ZN(n3469) );
  inv0d0 U351 ( .I(n5477), .ZN(n3318) );
  inv0d0 U352 ( .I(n7485), .ZN(n4369) );
  inv0d0 U353 ( .I(n8026), .ZN(n2907) );
  inv0d0 U354 ( .I(n7754), .ZN(n3532) );
  nd02d1 U355 ( .A1(n3411), .A2(n3413), .ZN(n5438) );
  nd02d1 U356 ( .A1(n4068), .A2(n4112), .ZN(n7573) );
  nd02d1 U357 ( .A1(n3005), .A2(n11858), .ZN(n4800) );
  inv0d0 U358 ( .I(n7123), .ZN(n3401) );
  inv0d0 U359 ( .I(n6215), .ZN(n3372) );
  inv0d0 U360 ( .I(n4872), .ZN(n2870) );
  inv0d0 U361 ( .I(n5031), .ZN(n4063) );
  inv0d0 U362 ( .I(n9523), .ZN(n2994) );
  inv0d0 U363 ( .I(n6391), .ZN(n3189) );
  inv0d0 U364 ( .I(n10643), .ZN(n3929) );
  inv0d0 U365 ( .I(n9235), .ZN(n3789) );
  inv0d0 U366 ( .I(n8112), .ZN(n4154) );
  buffd1 U367 ( .I(n690), .Z(n563) );
  buffd1 U368 ( .I(n690), .Z(n564) );
  buffd1 U369 ( .I(n690), .Z(n565) );
  buffd1 U370 ( .I(n689), .Z(n566) );
  buffd1 U371 ( .I(n689), .Z(n567) );
  buffd1 U372 ( .I(n689), .Z(n568) );
  buffd1 U373 ( .I(n688), .Z(n569) );
  buffd1 U374 ( .I(n688), .Z(n570) );
  buffd1 U375 ( .I(n688), .Z(n571) );
  buffd1 U376 ( .I(n687), .Z(n572) );
  buffd1 U377 ( .I(n687), .Z(n573) );
  buffd1 U378 ( .I(n694), .Z(n551) );
  buffd1 U379 ( .I(n694), .Z(n552) );
  buffd1 U380 ( .I(n694), .Z(n553) );
  buffd1 U381 ( .I(n693), .Z(n554) );
  buffd1 U382 ( .I(n693), .Z(n555) );
  buffd1 U383 ( .I(n693), .Z(n556) );
  buffd1 U384 ( .I(n692), .Z(n557) );
  buffd1 U385 ( .I(n692), .Z(n558) );
  buffd1 U386 ( .I(n692), .Z(n559) );
  buffd1 U387 ( .I(n691), .Z(n560) );
  buffd1 U388 ( .I(n691), .Z(n561) );
  buffd1 U389 ( .I(n691), .Z(n562) );
  buffd1 U390 ( .I(n682), .Z(n587) );
  buffd1 U391 ( .I(n682), .Z(n588) );
  buffd1 U392 ( .I(n682), .Z(n589) );
  buffd1 U393 ( .I(n681), .Z(n590) );
  buffd1 U394 ( .I(n681), .Z(n591) );
  buffd1 U395 ( .I(n680), .Z(n593) );
  buffd1 U396 ( .I(n680), .Z(n594) );
  buffd1 U397 ( .I(n680), .Z(n595) );
  buffd1 U398 ( .I(n679), .Z(n596) );
  buffd1 U399 ( .I(n679), .Z(n597) );
  buffd1 U400 ( .I(n686), .Z(n575) );
  buffd1 U401 ( .I(n686), .Z(n576) );
  buffd1 U402 ( .I(n686), .Z(n577) );
  buffd1 U403 ( .I(n685), .Z(n578) );
  buffd1 U404 ( .I(n685), .Z(n579) );
  buffd1 U405 ( .I(n685), .Z(n580) );
  buffd1 U406 ( .I(n684), .Z(n581) );
  buffd1 U407 ( .I(n684), .Z(n582) );
  buffd1 U408 ( .I(n683), .Z(n584) );
  buffd1 U409 ( .I(n683), .Z(n585) );
  buffd1 U410 ( .I(n683), .Z(n586) );
  buffd1 U411 ( .I(n687), .Z(n574) );
  buffd1 U412 ( .I(n681), .Z(n592) );
  buffd1 U413 ( .I(n679), .Z(n598) );
  buffd1 U414 ( .I(n665), .Z(n640) );
  buffd1 U415 ( .I(n665), .Z(n639) );
  buffd1 U416 ( .I(n665), .Z(n638) );
  buffd1 U417 ( .I(n666), .Z(n637) );
  buffd1 U418 ( .I(n666), .Z(n636) );
  buffd1 U419 ( .I(n666), .Z(n635) );
  buffd1 U420 ( .I(n667), .Z(n633) );
  buffd1 U421 ( .I(n667), .Z(n632) );
  buffd1 U422 ( .I(n668), .Z(n631) );
  buffd1 U423 ( .I(n668), .Z(n630) );
  buffd1 U424 ( .I(n668), .Z(n629) );
  buffd1 U425 ( .I(n669), .Z(n628) );
  buffd1 U426 ( .I(n667), .Z(n634) );
  buffd1 U427 ( .I(n662), .Z(n649) );
  buffd1 U428 ( .I(n661), .Z(n650) );
  buffd1 U429 ( .I(n661), .Z(n651) );
  buffd1 U430 ( .I(n660), .Z(n653) );
  buffd1 U431 ( .I(n660), .Z(n654) );
  buffd1 U432 ( .I(n660), .Z(n655) );
  buffd1 U433 ( .I(n662), .Z(n648) );
  buffd1 U434 ( .I(n662), .Z(n647) );
  buffd1 U435 ( .I(n663), .Z(n646) );
  buffd1 U436 ( .I(n663), .Z(n645) );
  buffd1 U437 ( .I(n663), .Z(n644) );
  buffd1 U438 ( .I(n664), .Z(n643) );
  buffd1 U439 ( .I(n664), .Z(n642) );
  buffd1 U440 ( .I(n664), .Z(n641) );
  buffd1 U441 ( .I(n661), .Z(n652) );
  buffd1 U442 ( .I(n674), .Z(n611) );
  buffd1 U443 ( .I(n675), .Z(n610) );
  buffd1 U444 ( .I(n675), .Z(n609) );
  buffd1 U445 ( .I(n675), .Z(n608) );
  buffd1 U446 ( .I(n676), .Z(n607) );
  buffd1 U447 ( .I(n676), .Z(n606) );
  buffd1 U448 ( .I(n678), .Z(n599) );
  buffd1 U449 ( .I(n678), .Z(n600) );
  buffd1 U450 ( .I(n678), .Z(n601) );
  buffd1 U451 ( .I(n677), .Z(n602) );
  buffd1 U452 ( .I(n677), .Z(n603) );
  buffd1 U453 ( .I(n677), .Z(n604) );
  buffd1 U454 ( .I(n676), .Z(n605) );
  buffd1 U455 ( .I(n669), .Z(n626) );
  buffd1 U456 ( .I(n670), .Z(n625) );
  buffd1 U457 ( .I(n670), .Z(n624) );
  buffd1 U458 ( .I(n670), .Z(n623) );
  buffd1 U459 ( .I(n671), .Z(n622) );
  buffd1 U460 ( .I(n671), .Z(n621) );
  buffd1 U461 ( .I(n672), .Z(n619) );
  buffd1 U462 ( .I(n672), .Z(n618) );
  buffd1 U463 ( .I(n672), .Z(n617) );
  buffd1 U464 ( .I(n673), .Z(n616) );
  buffd1 U465 ( .I(n673), .Z(n615) );
  buffd1 U466 ( .I(n673), .Z(n614) );
  buffd1 U467 ( .I(n674), .Z(n613) );
  buffd1 U468 ( .I(n674), .Z(n612) );
  buffd1 U469 ( .I(n671), .Z(n620) );
  buffd1 U470 ( .I(n669), .Z(n627) );
  inv0d0 U471 ( .I(n10613), .ZN(n4027) );
  inv0d0 U472 ( .I(n11037), .ZN(n3074) );
  inv0d0 U473 ( .I(n7197), .ZN(n3300) );
  nd02d1 U474 ( .A1(n3800), .A2(n9957), .ZN(n4417) );
  inv0d0 U475 ( .I(n5659), .ZN(n2960) );
  inv0d0 U476 ( .I(n9632), .ZN(n3934) );
  inv0d0 U477 ( .I(n8178), .ZN(n4281) );
  buffd1 U478 ( .I(n684), .Z(n583) );
  inv0d0 U479 ( .I(n4933), .ZN(n2981) );
  inv0d0 U480 ( .I(n7796), .ZN(n3451) );
  inv0d0 U481 ( .I(n7346), .ZN(n2851) );
  inv0d0 U482 ( .I(n8842), .ZN(n3294) );
  inv0d0 U483 ( .I(n6031), .ZN(n3837) );
  inv0d0 U484 ( .I(n9194), .ZN(n3740) );
  inv0d0 U485 ( .I(n11003), .ZN(n3214) );
  inv0d0 U486 ( .I(n10593), .ZN(n4013) );
  inv0d0 U487 ( .I(n4648), .ZN(n3173) );
  inv0d0 U488 ( .I(n6372), .ZN(n3177) );
  inv0d0 U489 ( .I(n7866), .ZN(n3290) );
  inv0d0 U490 ( .I(n6883), .ZN(n3915) );
  inv0d0 U491 ( .I(n10343), .ZN(n2897) );
  inv0d0 U492 ( .I(n11918), .ZN(n2875) );
  inv0d0 U493 ( .I(n11242), .ZN(n3449) );
  inv0d0 U494 ( .I(n5793), .ZN(n4195) );
  inv0d0 U495 ( .I(n4849), .ZN(n2931) );
  inv0d0 U496 ( .I(n7044), .ZN(n3553) );
  inv0d0 U497 ( .I(n7287), .ZN(n3082) );
  inv0d0 U498 ( .I(n4536), .ZN(n3365) );
  inv0d0 U499 ( .I(n6643), .ZN(n4026) );
  inv0d0 U500 ( .I(n9268), .ZN(n3554) );
  inv0d0 U501 ( .I(n6943), .ZN(n3841) );
  inv0d0 U502 ( .I(n7274), .ZN(n3057) );
  inv0d0 U503 ( .I(n6262), .ZN(n3394) );
  inv0d0 U504 ( .I(n5995), .ZN(n3935) );
  inv0d0 U505 ( .I(n11300), .ZN(n4789) );
  inv0d0 U506 ( .I(n11136), .ZN(n2860) );
  inv0d0 U507 ( .I(n8416), .ZN(n3867) );
  inv0d0 U508 ( .I(n4589), .ZN(n3320) );
  inv0d0 U509 ( .I(n7764), .ZN(n3562) );
  inv0d0 U510 ( .I(n9661), .ZN(n4793) );
  inv0d0 U511 ( .I(n10235), .ZN(n2947) );
  inv0d0 U512 ( .I(n7008), .ZN(n3653) );
  inv0d0 U513 ( .I(n8502), .ZN(n3476) );
  inv0d0 U514 ( .I(n6569), .ZN(n3069) );
  inv0d0 U515 ( .I(N5116), .ZN(n1397) );
  inv0d0 U516 ( .I(n5668), .ZN(n2971) );
  inv0d0 U517 ( .I(n7786), .ZN(n3432) );
  inv0d0 U518 ( .I(n7609), .ZN(n4002) );
  inv0d0 U519 ( .I(n6464), .ZN(n3052) );
  inv0d0 U520 ( .I(n6436), .ZN(n3042) );
  inv0d0 U521 ( .I(n7846), .ZN(n3386) );
  inv0d0 U522 ( .I(N5117), .ZN(n1398) );
  inv0d0 U523 ( .I(n11368), .ZN(n4253) );
  inv0d0 U524 ( .I(n11557), .ZN(n3886) );
  inv0d0 U525 ( .I(n8194), .ZN(n4247) );
  inv0d0 U526 ( .I(N5118), .ZN(n1399) );
  inv0d0 U527 ( .I(n5772), .ZN(n3955) );
  inv0d0 U528 ( .I(n11729), .ZN(n3385) );
  inv0d0 U529 ( .I(n4823), .ZN(n2932) );
  inv0d0 U530 ( .I(n8332), .ZN(n4036) );
  inv0d0 U531 ( .I(n6535), .ZN(n2920) );
  inv0d0 U532 ( .I(n10081), .ZN(n3396) );
  inv0d0 U533 ( .I(n7490), .ZN(n4368) );
  inv0d0 U534 ( .I(n4479), .ZN(n3423) );
  inv0d0 U535 ( .I(n8190), .ZN(n4274) );
  inv0d0 U536 ( .I(n6584), .ZN(n3228) );
  inv0d0 U537 ( .I(n10124), .ZN(n3172) );
  inv0d0 U538 ( .I(n9247), .ZN(n3535) );
  inv0d0 U539 ( .I(n5018), .ZN(n4186) );
  inv0d0 U540 ( .I(N5120), .ZN(n1400) );
  inv0d0 U541 ( .I(n1379), .ZN(N5120) );
  inv0d0 U542 ( .I(n5703), .ZN(n3071) );
  inv0d0 U543 ( .I(n7493), .ZN(n4280) );
  inv0d0 U544 ( .I(n6625), .ZN(n3830) );
  inv0d0 U545 ( .I(n10071), .ZN(n3407) );
  inv0d0 U546 ( .I(n7527), .ZN(n4146) );
  inv0d0 U547 ( .I(n8391), .ZN(n3833) );
  inv0d0 U548 ( .I(n5635), .ZN(n2924) );
  inv0d0 U549 ( .I(n5799), .ZN(n4215) );
  inv0d0 U550 ( .I(n4425), .ZN(n3725) );
  nd02d1 U551 ( .A1(n31), .A2(n512), .ZN(n10) );
  nd02d1 U552 ( .A1(n3647), .A2(n3648), .ZN(n3617) );
  buffd1 U553 ( .I(n391), .Z(n428) );
  buffd1 U554 ( .I(n391), .Z(n427) );
  buffd1 U555 ( .I(n391), .Z(n429) );
  buffd1 U556 ( .I(n392), .Z(n437) );
  buffd1 U557 ( .I(n393), .Z(n447) );
  buffd1 U558 ( .I(n393), .Z(n446) );
  buffd1 U559 ( .I(n392), .Z(n438) );
  buffd1 U560 ( .I(n393), .Z(n448) );
  buffd1 U561 ( .I(n394), .Z(n456) );
  buffd1 U562 ( .I(n394), .Z(n457) );
  buffd1 U563 ( .I(n3585), .Z(n950) );
  buffd1 U564 ( .I(n3585), .Z(n951) );
  buffd1 U565 ( .I(n3585), .Z(n949) );
  buffd1 U566 ( .I(n3584), .Z(n954) );
  buffd1 U567 ( .I(n3584), .Z(n952) );
  buffd1 U568 ( .I(n3584), .Z(n953) );
  inv0d0 U569 ( .I(N5285), .ZN(n2774) );
  nr02d1 U570 ( .A1(n505), .A2(n503), .ZN(n383) );
  inv0d0 U571 ( .I(n2713), .ZN(n2722) );
  buffd1 U572 ( .I(n838), .Z(n843) );
  buffd1 U573 ( .I(n838), .Z(n842) );
  buffd1 U574 ( .I(n838), .Z(n841) );
  buffd1 U575 ( .I(n839), .Z(n844) );
  buffd1 U576 ( .I(n4343), .Z(n826) );
  buffd1 U577 ( .I(n4343), .Z(n825) );
  buffd1 U578 ( .I(n4343), .Z(n824) );
  buffd1 U579 ( .I(n4258), .Z(n870) );
  buffd1 U580 ( .I(n4343), .Z(n827) );
  buffd1 U581 ( .I(n744), .Z(n749) );
  buffd1 U582 ( .I(n744), .Z(n748) );
  buffd1 U583 ( .I(n744), .Z(n747) );
  buffd1 U584 ( .I(n745), .Z(n750) );
  buffd1 U585 ( .I(n4258), .Z(n871) );
  buffd1 U586 ( .I(n4371), .Z(n720) );
  buffd1 U587 ( .I(n4371), .Z(n719) );
  buffd1 U588 ( .I(n4371), .Z(n718) );
  buffd1 U589 ( .I(n4371), .Z(n721) );
  buffd1 U590 ( .I(n4258), .Z(n872) );
  buffd1 U591 ( .I(n839), .Z(n846) );
  buffd1 U592 ( .I(n839), .Z(n845) );
  buffd1 U593 ( .I(n4354), .Z(n805) );
  buffd1 U594 ( .I(n4354), .Z(n804) );
  buffd1 U595 ( .I(n4354), .Z(n803) );
  buffd1 U596 ( .I(n4354), .Z(n806) );
  buffd1 U597 ( .I(n4343), .Z(n829) );
  buffd1 U598 ( .I(n4343), .Z(n828) );
  buffd1 U599 ( .I(n4343), .Z(n830) );
  buffd1 U600 ( .I(n745), .Z(n752) );
  buffd1 U601 ( .I(n745), .Z(n751) );
  buffd1 U602 ( .I(n780), .Z(n786) );
  buffd1 U603 ( .I(n780), .Z(n787) );
  buffd1 U604 ( .I(n779), .Z(n782) );
  buffd1 U605 ( .I(n779), .Z(n783) );
  buffd1 U606 ( .I(n779), .Z(n784) );
  buffd1 U607 ( .I(n780), .Z(n785) );
  buffd1 U608 ( .I(n4371), .Z(n723) );
  buffd1 U609 ( .I(n4371), .Z(n722) );
  buffd1 U610 ( .I(n781), .Z(n788) );
  buffd1 U611 ( .I(n4371), .Z(n724) );
  buffd1 U612 ( .I(n4354), .Z(n808) );
  buffd1 U613 ( .I(n4354), .Z(n807) );
  buffd1 U614 ( .I(n4354), .Z(n809) );
  inv0d0 U615 ( .I(n494), .ZN(n493) );
  inv0d0 U616 ( .I(reorder_start), .ZN(n494) );
  inv0d0 U617 ( .I(n3590), .ZN(n2753) );
  inv0d0 U618 ( .I(n3667), .ZN(n2759) );
  inv0d0 U619 ( .I(N4010), .ZN(N5108) );
  inv0d0 U620 ( .I(n1617), .ZN(n1620) );
  nr02d1 U621 ( .A1(n11966), .A2(n9538), .ZN(n4933) );
  nr02d1 U622 ( .A1(n7336), .A2(n3002), .ZN(n4810) );
  nr02d1 U623 ( .A1(n11229), .A2(n11231), .ZN(n6316) );
  nr02d1 U624 ( .A1(n6499), .A2(n11071), .ZN(n5619) );
  nr02d1 U625 ( .A1(n11056), .A2(n11053), .ZN(n9599) );
  nr02d1 U626 ( .A1(n8688), .A2(n6577), .ZN(n4721) );
  nr02d1 U627 ( .A1(n5050), .A2(n11277), .ZN(n4391) );
  nd12d1 U628 ( .A1(n11738), .A2(n11737), .ZN(n4586) );
  nr02d1 U629 ( .A1(n7335), .A2(n2844), .ZN(n5678) );
  nr02d1 U630 ( .A1(n9860), .A2(n5131), .ZN(n6883) );
  nr02d1 U631 ( .A1(n10327), .A2(n11155), .ZN(n8026) );
  nd03d1 U632 ( .A1(n3947), .A2(n4420), .A3(n4032), .ZN(n4415) );
  nr02d1 U633 ( .A1(n10279), .A2(n10280), .ZN(n8787) );
  nr02d1 U634 ( .A1(n8722), .A2(n6480), .ZN(n4764) );
  nd02d1 U635 ( .A1(n7972), .A2(n7973), .ZN(n7971) );
  nr02d1 U636 ( .A1(n3047), .A2(n6448), .ZN(n4715) );
  inv0d0 U637 ( .I(n4928), .ZN(n2827) );
  nr02d1 U638 ( .A1(n8919), .A2(n8909), .ZN(n6681) );
  nr02d1 U639 ( .A1(n6197), .A2(n6198), .ZN(n4528) );
  nr02d1 U640 ( .A1(n8731), .A2(n4778), .ZN(n6500) );
  nd02d1 U641 ( .A1(n7889), .A2(n3191), .ZN(n6391) );
  nr02d1 U642 ( .A1(n4586), .A2(n7163), .ZN(n6292) );
  nd02d1 U643 ( .A1(N14018), .A2(n3224), .ZN(n6588) );
  nr02d1 U644 ( .A1(n2852), .A2(n2912), .ZN(n9554) );
  nr02d1 U645 ( .A1(n9777), .A2(n11283), .ZN(n8104) );
  nr02d1 U646 ( .A1(n8943), .A2(n11348), .ZN(n6691) );
  nd02d1 U647 ( .A1(N14546), .A2(n3101), .ZN(n11071) );
  nr02d1 U648 ( .A1(n5477), .A2(n7386), .ZN(n6295) );
  nr02d1 U649 ( .A1(n10102), .A2(n10097), .ZN(n5487) );
  nr02d1 U650 ( .A1(n5027), .A2(n4061), .ZN(n8105) );
  nr02d1 U651 ( .A1(n4839), .A2(n2974), .ZN(n4838) );
  nd02d1 U652 ( .A1(n8839), .A2(n3297), .ZN(n8842) );
  nr02d1 U653 ( .A1(n6448), .A2(n8688), .ZN(n8683) );
  nr02d1 U654 ( .A1(n4778), .A2(n3014), .ZN(n4777) );
  nr02d1 U655 ( .A1(n4177), .A2(n5848), .ZN(n5023) );
  nd02d1 U656 ( .A1(N14850), .A2(n3001), .ZN(n7336) );
  nr02d1 U657 ( .A1(n8661), .A2(n6588), .ZN(n11003) );
  nr02d1 U658 ( .A1(n3732), .A2(n5279), .ZN(n6063) );
  nd12d1 U659 ( .A1(n1717), .A2(n3244), .ZN(n6372) );
  nd02d1 U660 ( .A1(n4721), .A2(n6448), .ZN(n4720) );
  nd02d1 U661 ( .A1(N15362), .A2(n2910), .ZN(n9562) );
  nd02d1 U662 ( .A1(N12418), .A2(n11679), .ZN(n8534) );
  nr02d1 U663 ( .A1(n4756), .A2(n10382), .ZN(n7287) );
  nd02d1 U664 ( .A1(n3419), .A2(n3366), .ZN(n4536) );
  nr02d1 U665 ( .A1(n6913), .A2(n5158), .ZN(n9632) );
  inv0d0 U666 ( .I(n2649), .ZN(N8246) );
  nd02d1 U667 ( .A1(n11137), .A2(n11190), .ZN(n4872) );
  nd12d1 U668 ( .A1(n2242), .A2(n9876), .ZN(n5995) );
  nd02d1 U669 ( .A1(N11196), .A2(n3808), .ZN(n9202) );
  nr02d1 U670 ( .A1(n8320), .A2(n5066), .ZN(n7614) );
  nd02d1 U671 ( .A1(n3562), .A2(n3538), .ZN(n6616) );
  nd02d1 U672 ( .A1(N11136), .A2(n3744), .ZN(n5287) );
  nr02d1 U673 ( .A1(n8059), .A2(n7898), .ZN(n4678) );
  nr02d1 U674 ( .A1(n11140), .A2(n11928), .ZN(n11918) );
  nd02d1 U675 ( .A1(n3373), .A2(n3411), .ZN(n6215) );
  nr02d1 U676 ( .A1(n9629), .A2(n10674), .ZN(n6031) );
  nd12d1 U677 ( .A1(n2545), .A2(n4201), .ZN(n5793) );
  nr02d1 U678 ( .A1(n5583), .A2(n4733), .ZN(n7274) );
  nd02d1 U679 ( .A1(n4065), .A2(n4064), .ZN(n5031) );
  nd02d1 U680 ( .A1(N14082), .A2(n3229), .ZN(n6584) );
  nd03d1 U681 ( .A1(n3560), .A2(n9998), .A3(n3537), .ZN(n4465) );
  nr02d1 U682 ( .A1(n11541), .A2(n4318), .ZN(n11550) );
  nd02d1 U683 ( .A1(n3301), .A2(n3302), .ZN(n7197) );
  inv0d0 U684 ( .I(n6460), .ZN(n3123) );
  nr02d1 U685 ( .A1(n6518), .A2(n6551), .ZN(n6521) );
  nr02d1 U686 ( .A1(n5316), .A2(n5750), .ZN(n5327) );
  nd02d1 U687 ( .A1(N11436), .A2(n3793), .ZN(n9227) );
  nr02d1 U688 ( .A1(n4499), .A2(n4995), .ZN(n4500) );
  nd02d1 U689 ( .A1(N15586), .A2(n2902), .ZN(n10343) );
  inv0d0 U690 ( .I(n7973), .ZN(n2927) );
  nr02d1 U691 ( .A1(n7313), .A2(n9512), .ZN(n4798) );
  nr02d1 U692 ( .A1(n11667), .A2(n4995), .ZN(n11669) );
  nr02d1 U693 ( .A1(n4849), .A2(n4932), .ZN(n4853) );
  inv0d0 U694 ( .I(n4850), .ZN(n2829) );
  nr02d1 U695 ( .A1(n7370), .A2(n6584), .ZN(n7259) );
  nd02d1 U696 ( .A1(n3319), .A2(n3321), .ZN(n5477) );
  nd02d1 U697 ( .A1(N14530), .A2(n10203), .ZN(n8722) );
  nd02d1 U698 ( .A1(n3402), .A2(n3404), .ZN(n7123) );
  nr02d1 U699 ( .A1(n11885), .A2(n4932), .ZN(n11896) );
  nd02d1 U700 ( .A1(n3406), .A2(n3408), .ZN(n5445) );
  nr02d1 U701 ( .A1(n5663), .A2(n4932), .ZN(n5674) );
  nd02d1 U702 ( .A1(n3066), .A2(n3123), .ZN(n6465) );
  nr02d1 U703 ( .A1(n7970), .A2(n7973), .ZN(n7300) );
  nd02d1 U704 ( .A1(n3868), .A2(n3869), .ZN(n8416) );
  nd02d1 U705 ( .A1(n3477), .A2(n5368), .ZN(n8502) );
  nr02d1 U706 ( .A1(n11869), .A2(n4998), .ZN(n11883) );
  nr02d1 U707 ( .A1(n5206), .A2(n9629), .ZN(n5211) );
  nd02d1 U708 ( .A1(N8096), .A2(n4832), .ZN(n9661) );
  nd02d1 U709 ( .A1(N12274), .A2(n3462), .ZN(n5402) );
  nd02d1 U710 ( .A1(n3065), .A2(n3122), .ZN(n4739) );
  nd02d1 U711 ( .A1(n3073), .A2(n10188), .ZN(n5703) );
  nr02d1 U712 ( .A1(n5649), .A2(n4998), .ZN(n5658) );
  nd02d1 U713 ( .A1(N8938), .A2(n4180), .ZN(n5831) );
  nd02d1 U714 ( .A1(n10788), .A2(n3545), .ZN(n5374) );
  nd02d1 U715 ( .A1(n3074), .A2(n3122), .ZN(n6569) );
  nd02d1 U716 ( .A1(n3843), .A2(n3844), .ZN(n6943) );
  nd02d1 U717 ( .A1(N11698), .A2(n3534), .ZN(n7754) );
  nd02d1 U718 ( .A1(n3388), .A2(n3393), .ZN(n7139) );
  nr02d1 U719 ( .A1(n9528), .A2(n2986), .ZN(n7326) );
  nr02d1 U720 ( .A1(n10734), .A2(n10735), .ZN(n9957) );
  nr02d1 U721 ( .A1(n6577), .A2(n4713), .ZN(n6436) );
  nd02d1 U722 ( .A1(N15058), .A2(n2980), .ZN(n7331) );
  nd03d1 U723 ( .A1(n3452), .A2(n3456), .A3(n3454), .ZN(n7796) );
  nr02d1 U724 ( .A1(n6996), .A2(n5750), .ZN(n7008) );
  nd02d1 U725 ( .A1(n2903), .A2(n2891), .ZN(n4891) );
  nr02d1 U726 ( .A1(n5374), .A2(n5366), .ZN(n4466) );
  nr02d1 U727 ( .A1(n4803), .A2(n7313), .ZN(n10235) );
  nr02d1 U728 ( .A1(n7211), .A2(n9607), .ZN(n8844) );
  nr02d1 U729 ( .A1(n6913), .A2(n11540), .ZN(n5161) );
  nd02d1 U730 ( .A1(N10536), .A2(n3960), .ZN(n8380) );
  nr02d1 U731 ( .A1(n8125), .A2(n6671), .ZN(n7493) );
  nr02d1 U732 ( .A1(n5006), .A2(n5015), .ZN(n7609) );
  nr02d1 U733 ( .A1(n9369), .A2(n11729), .ZN(n7846) );
  nr02d1 U734 ( .A1(n3245), .A2(n3244), .ZN(n4641) );
  nr02d1 U735 ( .A1(n6347), .A2(n7197), .ZN(n6342) );
  nr02d1 U736 ( .A1(n6480), .A2(n3108), .ZN(n6485) );
  nd02d1 U737 ( .A1(n5341), .A2(n4760), .ZN(n4765) );
  nr02d1 U738 ( .A1(n10067), .A2(n3408), .ZN(n10071) );
  nd02d1 U739 ( .A1(N12482), .A2(n6193), .ZN(n11242) );
  inv0d0 U740 ( .I(n6365), .ZN(n3250) );
  inv0d0 U741 ( .I(n5037), .ZN(n4165) );
  nd02d1 U742 ( .A1(n2829), .A2(n10280), .ZN(n4857) );
  nd02d1 U743 ( .A1(n7987), .A2(n4933), .ZN(n5668) );
  nr02d1 U744 ( .A1(n3451), .A2(n7792), .ZN(n4515) );
  nr02d1 U745 ( .A1(n8502), .A2(n3551), .ZN(n4476) );
  nd02d1 U746 ( .A1(N10716), .A2(n3879), .ZN(n10674) );
  nd02d1 U747 ( .A1(n3433), .A2(n3460), .ZN(n5404) );
  inv0d0 U748 ( .I(n9512), .ZN(n3005) );
  nd02d1 U749 ( .A1(n3387), .A2(n3395), .ZN(n11729) );
  nd02d1 U750 ( .A1(N12018), .A2(n3556), .ZN(n9268) );
  nr02d1 U751 ( .A1(n6286), .A2(n4978), .ZN(n6302) );
  nd03d1 U752 ( .A1(n4098), .A2(n8876), .A3(n4097), .ZN(n5040) );
  nd02d1 U753 ( .A1(N11810), .A2(n3563), .ZN(n7764) );
  nr02d1 U754 ( .A1(n4657), .A2(n5142), .ZN(n4669) );
  nd03d1 U755 ( .A1(n3742), .A2(n3809), .A3(n6073), .ZN(n9194) );
  nd02d1 U756 ( .A1(n4053), .A2(n11275), .ZN(n6643) );
  nr02d1 U757 ( .A1(n2875), .A2(n11186), .ZN(n8807) );
  nr02d1 U758 ( .A1(n8606), .A2(n5512), .ZN(n10942) );
  inv0d0 U759 ( .I(n5666), .ZN(n2970) );
  inv0d0 U760 ( .I(n5552), .ZN(n3224) );
  inv0d0 U761 ( .I(n7163), .ZN(n3323) );
  nr02d1 U762 ( .A1(n3024), .A2(n4697), .ZN(n4701) );
  nr02d1 U763 ( .A1(n7337), .A2(n9554), .ZN(n4860) );
  inv0d0 U764 ( .I(n10732), .ZN(n3800) );
  inv0d0 U765 ( .I(n4904), .ZN(n2888) );
  nr02d1 U766 ( .A1(n11792), .A2(n5142), .ZN(n11795) );
  nr02d1 U767 ( .A1(n7912), .A2(n3024), .ZN(n7914) );
  inv0d0 U768 ( .I(n4446), .ZN(n3530) );
  nd02d1 U769 ( .A1(N8910), .A2(n4181), .ZN(n8112) );
  nr02d1 U770 ( .A1(n7236), .A2(n6391), .ZN(n6386) );
  nd03d1 U771 ( .A1(n3569), .A2(n3530), .A3(n7027), .ZN(n7410) );
  nd02d1 U772 ( .A1(n10189), .A2(n3121), .ZN(n7950) );
  nd02d1 U773 ( .A1(n3368), .A2(n3418), .ZN(n6203) );
  nd02d1 U774 ( .A1(N8458), .A2(n8188), .ZN(n8190) );
  inv0d0 U775 ( .I(n2603), .ZN(n2606) );
  nd03d1 U776 ( .A1(n3880), .A2(n3879), .A3(n3834), .ZN(n8391) );
  nd02d1 U777 ( .A1(n3556), .A2(n3553), .ZN(n5371) );
  nd02d1 U778 ( .A1(n4264), .A2(n8991), .ZN(n5799) );
  nd02d1 U779 ( .A1(n3397), .A2(n3398), .ZN(n10081) );
  nd02d1 U780 ( .A1(n2925), .A2(n4786), .ZN(n5635) );
  inv0d0 U781 ( .I(n7539), .ZN(n4180) );
  inv0d0 U782 ( .I(n11409), .ZN(n4179) );
  nr02d1 U783 ( .A1(n6588), .A2(n5552), .ZN(n8653) );
  nd02d1 U784 ( .A1(n3011), .A2(n2927), .ZN(n4779) );
  nd02d1 U785 ( .A1(N11286), .A2(n3804), .ZN(n10726) );
  inv0d0 U786 ( .I(n6016), .ZN(n3828) );
  nd02d1 U787 ( .A1(n8991), .A2(n11385), .ZN(n8115) );
  nd02d1 U788 ( .A1(n8383), .A2(n3956), .ZN(n5772) );
  nd02d1 U789 ( .A1(N12194), .A2(n7064), .ZN(n7059) );
  inv0d0 U790 ( .I(n1951), .ZN(n1952) );
  inv0d0 U791 ( .I(n6406), .ZN(n3232) );
  nd02d1 U792 ( .A1(n11550), .A2(n7423), .ZN(n11557) );
  inv0d0 U793 ( .I(n8297), .ZN(n4108) );
  nd02d1 U794 ( .A1(n9277), .A2(n3424), .ZN(n4479) );
  nd02d1 U795 ( .A1(N8294), .A2(n4383), .ZN(n8171) );
  nr02d1 U796 ( .A1(n4579), .A2(n3391), .ZN(n7142) );
  nr02d1 U797 ( .A1(n9468), .A2(n6459), .ZN(n10181) );
  nd02d1 U798 ( .A1(n3414), .A2(n3416), .ZN(n4545) );
  nd02d1 U799 ( .A1(n2850), .A2(n8802), .ZN(n7340) );
  nd02d1 U800 ( .A1(n4810), .A2(n2998), .ZN(n8765) );
  inv0d0 U801 ( .I(n10097), .ZN(n3286) );
  nd02d1 U802 ( .A1(n6063), .A2(n6062), .ZN(n4425) );
  inv0d0 U803 ( .I(n10728), .ZN(n3802) );
  nd02d1 U804 ( .A1(N12002), .A2(n10795), .ZN(n7044) );
  nd02d1 U805 ( .A1(n4187), .A2(n4189), .ZN(n5018) );
  nd02d1 U806 ( .A1(n3863), .A2(n3865), .ZN(n9185) );
  nd02d1 U807 ( .A1(n3244), .A2(n7216), .ZN(n4648) );
  nd02d1 U808 ( .A1(n3291), .A2(n10935), .ZN(n7866) );
  nd02d1 U809 ( .A1(n4187), .A2(n10423), .ZN(n5810) );
  nr02d1 U810 ( .A1(n6372), .A2(n8620), .ZN(n9421) );
  inv0d0 U811 ( .I(n7337), .ZN(n2913) );
  inv0d0 U812 ( .I(n8651), .ZN(n3211) );
  inv0d0 U813 ( .I(n10382), .ZN(n3117) );
  inv0d0 U814 ( .I(n11189), .ZN(n2871) );
  nr02d1 U815 ( .A1(n5383), .A2(n5388), .ZN(n8509) );
  inv0d0 U816 ( .I(n5562), .ZN(n3231) );
  nr02d1 U817 ( .A1(n9565), .A2(n8821), .ZN(n8006) );
  inv0d0 U818 ( .I(n7236), .ZN(n3241) );
  nd02d1 U819 ( .A1(n3227), .A2(n9453), .ZN(n6431) );
  nr02d1 U820 ( .A1(n10003), .A2(n9261), .ZN(n7035) );
  nr02d1 U821 ( .A1(n5317), .A2(n5319), .ZN(n6999) );
  inv0d0 U822 ( .I(n7211), .ZN(n3168) );
  inv0d0 U823 ( .I(n6557), .ZN(n3106) );
  inv0d0 U824 ( .I(n8021), .ZN(n2898) );
  nd02d1 U825 ( .A1(n3836), .A2(n3880), .ZN(n5206) );
  nd03d1 U826 ( .A1(n3472), .A2(n3474), .A3(n3473), .ZN(n5383) );
  inv0d0 U827 ( .I(n5418), .ZN(n3446) );
  nd12d1 U828 ( .A1(n11), .A2(n4269), .ZN(n11368) );
  nr04d1 U829 ( .A1(n1248), .A2(n2579), .A3(n1326), .A4(n1282), .ZN(n11) );
  nd02d1 U830 ( .A1(N14466), .A2(n3093), .ZN(n11056) );
  nr02d1 U831 ( .A1(n8547), .A2(n4536), .ZN(n8544) );
  inv0d0 U832 ( .I(n10280), .ZN(n2849) );
  inv0d0 U833 ( .I(n9438), .ZN(n3238) );
  nr02d1 U834 ( .A1(n4127), .A2(n4497), .ZN(n8296) );
  inv0d0 U835 ( .I(n12060), .ZN(n3957) );
  inv0d0 U836 ( .I(n10188), .ZN(n3121) );
  nr02d1 U837 ( .A1(n4423), .A2(n4605), .ZN(n4616) );
  inv0d0 U838 ( .I(n7569), .ZN(n4116) );
  nd02d1 U839 ( .A1(n3060), .A2(n6459), .ZN(n4731) );
  inv0d0 U840 ( .I(n10663), .ZN(n3956) );
  inv0d0 U841 ( .I(n7948), .ZN(n3054) );
  inv0d0 U842 ( .I(n11009), .ZN(n3227) );
  inv0d0 U843 ( .I(n5239), .ZN(n3873) );
  nd02d1 U844 ( .A1(n3409), .A2(n3410), .ZN(n10067) );
  inv0d0 U845 ( .I(n8337), .ZN(n4042) );
  nd02d1 U846 ( .A1(n11883), .A2(n4936), .ZN(n11885) );
  nd02d1 U847 ( .A1(n5658), .A2(n4936), .ZN(n5663) );
  inv0d0 U848 ( .I(n4778), .ZN(n3103) );
  nd02d1 U849 ( .A1(n11737), .A2(n11738), .ZN(n10090) );
  nr02d1 U850 ( .A1(n7357), .A2(n7358), .ZN(n4824) );
  inv0d0 U851 ( .I(n8507), .ZN(n3467) );
  inv0d0 U852 ( .I(n7963), .ZN(n3084) );
  nd03d1 U853 ( .A1(n3536), .A2(n7764), .A3(n3538), .ZN(n9247) );
  nd02d1 U854 ( .A1(n3394), .A2(n3398), .ZN(n7141) );
  nd02d1 U855 ( .A1(n10359), .A2(n2982), .ZN(n9543) );
  nd02d1 U856 ( .A1(n7877), .A2(n3243), .ZN(n7225) );
  nd03d1 U857 ( .A1(n3127), .A2(n3054), .A3(n3058), .ZN(n6464) );
  nd03d1 U858 ( .A1(n3290), .A2(n4623), .A3(n3284), .ZN(n4613) );
  inv0d0 U859 ( .I(n5027), .ZN(n4170) );
  nd02d1 U860 ( .A1(n3005), .A2(n7313), .ZN(n11858) );
  nd02d1 U861 ( .A1(n3367), .A2(n3416), .ZN(n7817) );
  inv0d0 U862 ( .I(n11672), .ZN(n3438) );
  nd02d1 U863 ( .A1(n11868), .A2(n4404), .ZN(n11869) );
  nd02d1 U864 ( .A1(n5646), .A2(n4404), .ZN(n5649) );
  nd02d1 U865 ( .A1(n11190), .A2(n2861), .ZN(n11136) );
  nd03d1 U866 ( .A1(n3175), .A2(n6377), .A3(n3173), .ZN(n10124) );
  nd02d1 U867 ( .A1(n4007), .A2(n9098), .ZN(n5055) );
  nd02d1 U868 ( .A1(n4029), .A2(n11275), .ZN(n10613) );
  inv0d0 U869 ( .I(n4795), .ZN(n2944) );
  nd02d1 U870 ( .A1(N9936), .A2(n4051), .ZN(n9836) );
  inv0d0 U871 ( .I(n11966), .ZN(n2980) );
  inv0d0 U872 ( .I(n8731), .ZN(n3105) );
  nd02d1 U873 ( .A1(n3035), .A2(n10161), .ZN(n4702) );
  inv0d0 U874 ( .I(n6059), .ZN(n3721) );
  inv0d0 U875 ( .I(n11954), .ZN(n2894) );
  inv0d0 U876 ( .I(n6478), .ZN(n3094) );
  inv0d0 U877 ( .I(n5951), .ZN(n3999) );
  inv0d0 U878 ( .I(n10910), .ZN(n3330) );
  nd02d1 U879 ( .A1(N9741), .A2(n4014), .ZN(n10593) );
  nd02d1 U880 ( .A1(n4404), .A2(n4805), .ZN(n4823) );
  nd02d1 U881 ( .A1(N14338), .A2(n3122), .ZN(n11037) );
  nd02d1 U882 ( .A1(n3321), .A2(n3323), .ZN(n4589) );
  nd02d1 U883 ( .A1(n5487), .A2(n3291), .ZN(n9394) );
  inv0d0 U884 ( .I(n7417), .ZN(n3856) );
  nd02d1 U885 ( .A1(n3097), .A2(n6499), .ZN(n4943) );
  nd02d1 U886 ( .A1(n3678), .A2(n3517), .ZN(n8460) );
  inv0d0 U887 ( .I(n6440), .ZN(n3035) );
  nd02d1 U888 ( .A1(n5541), .A2(n3205), .ZN(n4680) );
  inv0d0 U889 ( .I(n5512), .ZN(n3302) );
  nd02d1 U890 ( .A1(n4046), .A2(n10617), .ZN(n8332) );
  inv0d0 U891 ( .I(n10161), .ZN(n3037) );
  nd02d1 U892 ( .A1(n3240), .A2(n3205), .ZN(n11803) );
  nd02d1 U893 ( .A1(n8228), .A2(n4264), .ZN(n7527) );
  nd02d1 U894 ( .A1(n3433), .A2(n3434), .ZN(n7786) );
  nd02d1 U895 ( .A1(n11357), .A2(n4247), .ZN(n6710) );
  nd02d1 U896 ( .A1(n3435), .A2(n3459), .ZN(n9303) );
  inv0d0 U897 ( .I(n6237), .ZN(n3375) );
  inv0d0 U898 ( .I(n6314), .ZN(n3314) );
  inv0d0 U899 ( .I(n7581), .ZN(n4104) );
  inv0d0 U900 ( .I(n6416), .ZN(n3208) );
  inv0d0 U901 ( .I(n8016), .ZN(n2903) );
  inv0d0 U902 ( .I(n5416), .ZN(n3442) );
  nr02d1 U903 ( .A1(n6987), .A2(n4407), .ZN(n10716) );
  inv0d0 U904 ( .I(n4623), .ZN(n3293) );
  inv0d0 U905 ( .I(n6487), .ZN(n3111) );
  inv0d0 U906 ( .I(n4840), .ZN(n2983) );
  inv0d0 U907 ( .I(n7652), .ZN(n3964) );
  inv0d0 U908 ( .I(n11385), .ZN(n4201) );
  nd02d1 U909 ( .A1(n3419), .A2(n3364), .ZN(n5429) );
  nd02d1 U910 ( .A1(n3395), .A2(n3397), .ZN(n6262) );
  inv0d0 U911 ( .I(n8756), .ZN(n3004) );
  nd02d1 U912 ( .A1(n3790), .A2(n3789), .ZN(n11623) );
  nd02d1 U913 ( .A1(N10296), .A2(n3930), .ZN(n10643) );
  nd02d1 U914 ( .A1(N11241), .A2(n3764), .ZN(n9207) );
  inv0d0 U915 ( .I(n4935), .ZN(n2818) );
  nd02d1 U916 ( .A1(N8497), .A2(n4248), .ZN(n8194) );
  inv0d0 U917 ( .I(n4783), .ZN(n2925) );
  nd02d1 U918 ( .A1(n7259), .A2(n3229), .ZN(n9449) );
  nd02d1 U919 ( .A1(N8798), .A2(n4190), .ZN(n5805) );
  inv0d0 U920 ( .I(n5848), .ZN(n4176) );
  inv0d0 U921 ( .I(n6942), .ZN(n3832) );
  inv0d0 U922 ( .I(n9221), .ZN(n3798) );
  nd02d1 U923 ( .A1(n2998), .A2(n2995), .ZN(n9523) );
  nd02d1 U924 ( .A1(n3831), .A2(n3881), .ZN(n6625) );
  nd02d1 U925 ( .A1(n4373), .A2(n4369), .ZN(n7490) );
  nd02d1 U926 ( .A1(N11406), .A2(n3798), .ZN(n9222) );
  inv0d0 U927 ( .I(n5610), .ZN(n3087) );
  inv0d0 U928 ( .I(n7935), .ZN(n3060) );
  inv0d0 U929 ( .I(n7401), .ZN(n3434) );
  inv0d0 U930 ( .I(n10812), .ZN(n3474) );
  inv0d0 U931 ( .I(n6834), .ZN(n4098) );
  nd03d1 U932 ( .A1(n3323), .A2(n7857), .A3(n3321), .ZN(n7154) );
  inv0d0 U933 ( .I(n9437), .ZN(n3205) );
  inv0d0 U934 ( .I(n7890), .ZN(n3199) );
  nd02d1 U935 ( .A1(N8085), .A2(n4835), .ZN(n11300) );
  nd02d1 U936 ( .A1(n4149), .A2(n9008), .ZN(n10527) );
  inv0d0 U937 ( .I(n7428), .ZN(n3945) );
  inv0d0 U938 ( .I(n7987), .ZN(n2969) );
  nd02d1 U939 ( .A1(n3834), .A2(n5211), .ZN(n4402) );
  inv0d0 U940 ( .I(n8151), .ZN(n4604) );
  inv0d0 U941 ( .I(n6860), .ZN(n4054) );
  inv0d0 U942 ( .I(n8707), .ZN(n3076) );
  nd02d1 U943 ( .A1(n3178), .A2(n3177), .ZN(n8622) );
  inv0d0 U944 ( .I(n8526), .ZN(n3460) );
  inv0d0 U945 ( .I(n6122), .ZN(n3575) );
  inv0d0 U946 ( .I(n8672), .ZN(n3043) );
  aor211d1 U947 ( .C1(n1192), .C2(n1137), .A(n1280), .B(n1227), .Z(n12) );
  inv0d0 U948 ( .I(n8030), .ZN(n2940) );
  inv0d0 U949 ( .I(n11142), .ZN(n2910) );
  inv0d0 U950 ( .I(n10414), .ZN(n4033) );
  inv0d0 U951 ( .I(n4667), .ZN(n3188) );
  inv0d0 U952 ( .I(n8081), .ZN(n4692) );
  inv0d0 U953 ( .I(n6424), .ZN(n3222) );
  aor211d1 U954 ( .C1(n1192), .C2(n1138), .A(n1281), .B(n1256), .Z(n13) );
  inv0d0 U955 ( .I(n8893), .ZN(n4858) );
  inv0d0 U956 ( .I(n7357), .ZN(n2962) );
  inv0d0 U957 ( .I(n8821), .ZN(n2878) );
  inv0d0 U958 ( .I(n6515), .ZN(n2952) );
  inv0d0 U959 ( .I(n4863), .ZN(n2856) );
  inv0d0 U960 ( .I(n8241), .ZN(n4182) );
  inv0d0 U961 ( .I(n10734), .ZN(n3777) );
  inv0d0 U962 ( .I(n9687), .ZN(n4384) );
  nd02d1 U963 ( .A1(n8216), .A2(n4260), .ZN(n8964) );
  inv0d0 U964 ( .I(n10847), .ZN(n3443) );
  nd02d1 U965 ( .A1(n3405), .A2(n3409), .ZN(n6223) );
  inv0d1 U966 ( .I(n1315), .ZN(n1300) );
  inv0d1 U967 ( .I(n1215), .ZN(n1202) );
  inv0d0 U968 ( .I(n8344), .ZN(n4045) );
  inv0d1 U969 ( .I(n1316), .ZN(n1306) );
  inv0d1 U970 ( .I(n1169), .ZN(n1160) );
  inv0d1 U971 ( .I(n1259), .ZN(n1227) );
  inv0d1 U972 ( .I(n1310), .ZN(n1273) );
  inv0d1 U973 ( .I(n1211), .ZN(n1185) );
  inv0d0 U974 ( .I(n7386), .ZN(n3316) );
  nd02d1 U975 ( .A1(n3569), .A2(n3530), .ZN(n9243) );
  inv0d0 U976 ( .I(n9929), .ZN(n3865) );
  inv0d0 U977 ( .I(n10544), .ZN(n4175) );
  inv0d0 U978 ( .I(n10640), .ZN(n3933) );
  inv0d0 U979 ( .I(n10357), .ZN(n2982) );
  inv0d0 U980 ( .I(n6029), .ZN(n3881) );
  nd02d1 U981 ( .A1(n3782), .A2(n6111), .ZN(n7742) );
  inv0d0 U982 ( .I(n5326), .ZN(n3793) );
  inv0d0 U983 ( .I(n4409), .ZN(n3840) );
  inv0d0 U984 ( .I(n5115), .ZN(n3909) );
  inv0d0 U985 ( .I(n8320), .ZN(n4015) );
  inv0d0 U986 ( .I(n9336), .ZN(n3411) );
  inv0d0 U987 ( .I(n5087), .ZN(n4051) );
  inv0d0 U988 ( .I(n9472), .ZN(n3070) );
  inv0d0 U989 ( .I(n5004), .ZN(n4681) );
  inv0d0 U990 ( .I(n6987), .ZN(n3805) );
  inv0d0 U991 ( .I(n8031), .ZN(n2939) );
  inv0d0 U992 ( .I(n12042), .ZN(n3534) );
  inv0d0 U993 ( .I(n4995), .ZN(n4438) );
  inv0d0 U994 ( .I(n4508), .ZN(n3457) );
  inv0d0 U995 ( .I(n6527), .ZN(n2997) );
  inv0d0 U996 ( .I(n7857), .ZN(n3319) );
  inv0d0 U997 ( .I(n7358), .ZN(n2990) );
  inv0d0 U998 ( .I(n6634), .ZN(n5093) );
  inv0d0 U999 ( .I(n6118), .ZN(n3684) );
  inv0d0 U1000 ( .I(n4664), .ZN(n3183) );
  inv0d0 U1001 ( .I(n11137), .ZN(n2868) );
  inv0d0 U1002 ( .I(n4601), .ZN(n3313) );
  inv0d0 U1003 ( .I(n11039), .ZN(n3075) );
  nr02d1 U1004 ( .A1(n2796), .A2(n8707), .ZN(n8703) );
  inv0d0 U1005 ( .I(n5796), .ZN(n4231) );
  nd02d1 U1006 ( .A1(n3166), .A2(n3297), .ZN(n9410) );
  inv0d0 U1007 ( .I(n6197), .ZN(n3364) );
  inv0d0 U1008 ( .I(n10963), .ZN(n3248) );
  inv0d0 U1009 ( .I(n11873), .ZN(n2992) );
  inv0d0 U1010 ( .I(n7667), .ZN(n3943) );
  nd02d1 U1011 ( .A1(n6928), .A2(n7423), .ZN(n6940) );
  inv0d0 U1012 ( .I(n11126), .ZN(n2912) );
  inv0d0 U1013 ( .I(n6094), .ZN(n3773) );
  nd02d1 U1014 ( .A1(n3932), .A2(n3928), .ZN(n9872) );
  inv0d0 U1015 ( .I(n9896), .ZN(n3823) );
  inv0d0 U1016 ( .I(n5893), .ZN(n4124) );
  inv0d0 U1017 ( .I(n5305), .ZN(n3804) );
  inv0d0 U1018 ( .I(n5583), .ZN(n3056) );
  inv0d0 U1019 ( .I(n5050), .ZN(n4004) );
  inv0d0 U1020 ( .I(n5214), .ZN(n3844) );
  inv0d0 U1021 ( .I(n9402), .ZN(n3308) );
  inv0d0 U1022 ( .I(n9860), .ZN(n3914) );
  nd02d1 U1023 ( .A1(n3795), .A2(n3777), .ZN(n5328) );
  inv0d0 U1024 ( .I(n5017), .ZN(n4082) );
  inv0d0 U1025 ( .I(n5510), .ZN(n3165) );
  inv0d0 U1026 ( .I(n6786), .ZN(n4113) );
  inv0d0 U1027 ( .I(n4763), .ZN(n3089) );
  inv0d0 U1028 ( .I(n11140), .ZN(n2877) );
  nd02d1 U1029 ( .A1(n8131), .A2(n4835), .ZN(n8137) );
  inv0d0 U1030 ( .I(n4837), .ZN(n2968) );
  inv0d1 U1031 ( .I(n985), .ZN(n962) );
  inv0d0 U1032 ( .I(n5412), .ZN(n3459) );
  inv0d0 U1033 ( .I(n11853), .ZN(n2938) );
  inv0d0 U1034 ( .I(n8649), .ZN(n3207) );
  nd02d1 U1035 ( .A1(n3517), .A2(n3708), .ZN(n5349) );
  inv0d0 U1036 ( .I(n4534), .ZN(n3350) );
  inv0d0 U1037 ( .I(n12003), .ZN(n4426) );
  inv0d0 U1038 ( .I(n6950), .ZN(n3850) );
  inv0d0 U1039 ( .I(n9652), .ZN(n5314) );
  inv0d0 U1040 ( .I(n7277), .ZN(n3055) );
  inv0d0 U1041 ( .I(n8146), .ZN(n4816) );
  inv0d0 U1042 ( .I(n8616), .ZN(n3299) );
  inv0d0 U1045 ( .I(n6347), .ZN(n3298) );
  inv0d0 U1046 ( .I(n8464), .ZN(n3570) );
  inv0d0 U1047 ( .I(n5820), .ZN(n4747) );
  inv0d1 U1048 ( .I(n991), .ZN(n979) );
  inv0d1 U1049 ( .I(n985), .ZN(n963) );
  inv0d0 U1050 ( .I(n8008), .ZN(n2884) );
  inv0d0 U1051 ( .I(n9309), .ZN(n3452) );
  inv0d1 U1052 ( .I(n992), .ZN(n981) );
  inv0d1 U1053 ( .I(n991), .ZN(n980) );
  inv0d0 U1054 ( .I(n5319), .ZN(n3799) );
  inv0d0 U1055 ( .I(n4579), .ZN(n3271) );
  inv0d0 U1056 ( .I(n6542), .ZN(n2978) );
  inv0d0 U1057 ( .I(n5177), .ZN(n3950) );
  inv0d1 U1058 ( .I(n992), .ZN(n982) );
  inv0d0 U1061 ( .I(n5137), .ZN(n3920) );
  nd02d1 U1066 ( .A1(n7291), .A2(n5341), .ZN(n7303) );
  inv0d0 U1069 ( .I(n6377), .ZN(n3179) );
  inv0d0 U1072 ( .I(n6741), .ZN(n4214) );
  inv0d0 U1075 ( .I(n5020), .ZN(n4149) );
  inv0d0 U1078 ( .I(n9737), .ZN(n4196) );
  inv0d0 U1080 ( .I(n11791), .ZN(n3242) );
  inv0d0 U1081 ( .I(n9696), .ZN(n4279) );
  inv0d0 U1082 ( .I(n6551), .ZN(n4404) );
  inv0d1 U1083 ( .I(n989), .ZN(n973) );
  inv0d1 U1084 ( .I(n985), .ZN(n964) );
  inv0d0 U1085 ( .I(n1720), .ZN(N13682) );
  inv0d0 U1086 ( .I(n5244), .ZN(n3872) );
  inv0d1 U1087 ( .I(n987), .ZN(n969) );
  inv0d1 U1088 ( .I(n988), .ZN(n971) );
  inv0d1 U1089 ( .I(n988), .ZN(n972) );
  inv0d1 U1090 ( .I(n987), .ZN(n970) );
  inv0d1 U1093 ( .I(n989), .ZN(n974) );
  inv0d1 U1096 ( .I(n986), .ZN(n965) );
  inv0d1 U1099 ( .I(n986), .ZN(n966) );
  inv0d0 U1102 ( .I(n11053), .ZN(n3093) );
  inv0d0 U1105 ( .I(n5881), .ZN(n4064) );
  inv0d0 U1108 ( .I(n9468), .ZN(n3058) );
  inv0d1 U1111 ( .I(n986), .ZN(n967) );
  inv0d0 U1114 ( .I(n7362), .ZN(n3086) );
  inv0d0 U1117 ( .I(n7590), .ZN(n4085) );
  inv0d1 U1118 ( .I(n987), .ZN(n968) );
  inv0d0 U1119 ( .I(n5286), .ZN(n3809) );
  inv0d0 U1120 ( .I(n6739), .ZN(n4514) );
  inv0d0 U1122 ( .I(n10722), .ZN(n3764) );
  inv0d0 U1124 ( .I(n5153), .ZN(n3930) );
  inv0d0 U1125 ( .I(n9491), .ZN(n3014) );
  inv0d0 U1126 ( .I(n990), .ZN(n976) );
  inv0d0 U1128 ( .I(n11010), .ZN(n3030) );
  inv0d0 U1129 ( .I(n10322), .ZN(n2885) );
  inv0d0 U1131 ( .I(n990), .ZN(n975) );
  inv0d0 U1133 ( .I(n7653), .ZN(n3911) );
  inv0d0 U1135 ( .I(n11619), .ZN(n3787) );
  inv0d0 U1139 ( .I(n5032), .ZN(n4068) );
  inv0d0 U1153 ( .I(n7315), .ZN(n2956) );
  inv0d0 U1154 ( .I(n7216), .ZN(n3245) );
  inv0d0 U1155 ( .I(n7214), .ZN(n3163) );
  inv0d0 U1159 ( .I(n990), .ZN(n977) );
  inv0d0 U1160 ( .I(n5019), .ZN(n4112) );
  inv0d0 U1161 ( .I(n10661), .ZN(n3962) );
  inv0d0 U1162 ( .I(n8688), .ZN(n3051) );
  inv0d0 U1165 ( .I(n6564), .ZN(n3113) );
  inv0d0 U1167 ( .I(n5710), .ZN(n3201) );
  inv0d0 U1170 ( .I(n8597), .ZN(n3259) );
  inv0d0 U1171 ( .I(n6730), .ZN(n4261) );
  inv0d0 U1173 ( .I(n5363), .ZN(n3545) );
  inv0d0 U1174 ( .I(n5089), .ZN(n4481) );
  inv0d0 U1176 ( .I(n7522), .ZN(n4290) );
  inv0d0 U1177 ( .I(n11549), .ZN(n3952) );
  inv0d0 U1180 ( .I(n7031), .ZN(n3567) );
  inv0d0 U1191 ( .I(n9939), .ZN(n3808) );
  inv0d0 U1202 ( .I(n6754), .ZN(n4213) );
  inv0d0 U1203 ( .I(n5187), .ZN(n3819) );
  inv0d0 U1204 ( .I(n11484), .ZN(n4014) );
  inv0d0 U1242 ( .I(n8343), .ZN(n4038) );
  inv0d0 U1264 ( .I(n6791), .ZN(n4071) );
  inv0d0 U1280 ( .I(n5915), .ZN(n4079) );
  inv0d0 U1295 ( .I(n4740), .ZN(n3023) );
  inv0d0 U1312 ( .I(n6615), .ZN(n3560) );
  inv0d0 U1315 ( .I(n7972), .ZN(n2935) );
  inv0d0 U1328 ( .I(n10869), .ZN(n3414) );
  inv0d0 U1349 ( .I(n10350), .ZN(n2909) );
  inv0d0 U1350 ( .I(n991), .ZN(n978) );
  inv0d0 U1355 ( .I(n4615), .ZN(n3284) );
  inv0d0 U1372 ( .I(n4495), .ZN(n3468) );
  inv0d0 U1385 ( .I(n7309), .ZN(n2922) );
  inv0d0 U1418 ( .I(n10386), .ZN(n3045) );
  inv0d0 U1451 ( .I(n5368), .ZN(n3555) );
  inv0d0 U1458 ( .I(n5123), .ZN(n3913) );
  inv0d0 U1485 ( .I(n11541), .ZN(n3910) );
  inv0d0 U1518 ( .I(n9776), .ZN(n4118) );
  inv0d0 U1521 ( .I(n11439), .ZN(n4138) );
  inv0d0 U1534 ( .I(n9294), .ZN(n3464) );
  inv0d0 U1553 ( .I(n9791), .ZN(n4110) );
  inv0d0 U1586 ( .I(n7898), .ZN(n3202) );
  inv0d0 U1614 ( .I(n11348), .ZN(n4233) );
  inv0d0 U1616 ( .I(n6145), .ZN(n3557) );
  inv0d0 U1621 ( .I(n8383), .ZN(n3958) );
  inv0d0 U1622 ( .I(n8110), .ZN(n4166) );
  inv0d0 U1623 ( .I(n8043), .ZN(n2946) );
  inv0d0 U1630 ( .I(n7070), .ZN(n3489) );
  inv0d0 U1657 ( .I(n6480), .ZN(n3109) );
  inv0d0 U1660 ( .I(n6233), .ZN(n3359) );
  inv0d0 U1690 ( .I(n4602), .ZN(n3279) );
  inv0d0 U1692 ( .I(n8922), .ZN(n4365) );
  inv0d0 U1693 ( .I(n10327), .ZN(n2906) );
  inv0d0 U1694 ( .I(n5334), .ZN(n3785) );
  inv0d0 U1727 ( .I(n7631), .ZN(n4050) );
  inv0d0 U1728 ( .I(n7126), .ZN(n3354) );
  inv0d0 U1729 ( .I(n6727), .ZN(n4256) );
  inv0d0 U1730 ( .I(n7850), .ZN(n3274) );
  inv0d0 U1733 ( .I(n4467), .ZN(n4310) );
  inv0d0 U1735 ( .I(n11649), .ZN(n3508) );
  inv0d0 U1737 ( .I(n1761), .ZN(n1764) );
  inv0d0 U1739 ( .I(n1213), .ZN(n1209) );
  inv0d0 U1740 ( .I(n10339), .ZN(n2893) );
  inv0d0 U1742 ( .I(n11283), .ZN(n4168) );
  inv0d0 U1744 ( .I(n1437), .ZN(n1440) );
  inv0d0 U1746 ( .I(n8726), .ZN(n3102) );
  inv0d0 U1748 ( .I(n6757), .ZN(n4181) );
  inv0d0 U1750 ( .I(n9919), .ZN(n3851) );
  inv0d0 U1752 ( .I(n5127), .ZN(n3973) );
  inv0d0 U1754 ( .I(n5180), .ZN(n3960) );
  inv0d0 U1756 ( .I(n8094), .ZN(n4320) );
  inv0d0 U1757 ( .I(n11287), .ZN(n4160) );
  inv0d0 U1759 ( .I(n4981), .ZN(n5389) );
  inv0d0 U1761 ( .I(n6254), .ZN(n3383) );
  inv0d0 U1763 ( .I(n10463), .ZN(n4576) );
  inv0d0 U1764 ( .I(n4888), .ZN(n2883) );
  inv0d0 U1766 ( .I(n11231), .ZN(n3281) );
  inv0d0 U1768 ( .I(n9761), .ZN(n4173) );
  inv0d0 U1770 ( .I(n11579), .ZN(n3883) );
  inv0d0 U1772 ( .I(n6961), .ZN(n3869) );
  inv0d0 U1774 ( .I(n5395), .ZN(n3462) );
  nd02d1 U1776 ( .A1(n3834), .A2(n3832), .ZN(n9153) );
  inv0d0 U1778 ( .I(n4688), .ZN(n3158) );
  inv0d0 U1780 ( .I(n11693), .ZN(n3348) );
  inv0d0 U1782 ( .I(n5976), .ZN(n4043) );
  inv0d0 U1784 ( .I(n9839), .ZN(n4047) );
  inv0d0 U1786 ( .I(n6109), .ZN(n3782) );
  inv0d0 U1789 ( .I(n5699), .ZN(n5341) );
  inv0d0 U1792 ( .I(n5162), .ZN(n3971) );
  inv0d0 U1795 ( .I(n5007), .ZN(n4007) );
  inv0d0 U1798 ( .I(n10370), .ZN(n2948) );
  inv0d0 U1801 ( .I(n5492), .ZN(n3292) );
  inv0d0 U1802 ( .I(n7041), .ZN(n3542) );
  inv0d0 U1803 ( .I(n1262), .ZN(n1257) );
  inv0d0 U1804 ( .I(n11939), .ZN(n2834) );
  inv0d0 U1805 ( .I(n7650), .ZN(n3969) );
  inv0d0 U1807 ( .I(n5297), .ZN(n3759) );
  inv0d0 U1809 ( .I(n11366), .ZN(n4228) );
  inv0d0 U1810 ( .I(n10120), .ZN(n3166) );
  inv0d0 U1812 ( .I(n10912), .ZN(n3275) );
  inv0d0 U1813 ( .I(n11952), .ZN(n2900) );
  inv0d0 U1814 ( .I(n7905), .ZN(n3155) );
  inv0d0 U1815 ( .I(n6829), .ZN(n4091) );
  inv0d0 U1816 ( .I(n6022), .ZN(n3882) );
  inv0d0 U1826 ( .I(n6066), .ZN(n3734) );
  inv0d0 U1837 ( .I(n11540), .ZN(n3936) );
  inv0d0 U1838 ( .I(n9670), .ZN(n4568) );
  inv0d0 U1840 ( .I(n7700), .ZN(n3853) );
  inv0d0 U1842 ( .I(n8322), .ZN(n4018) );
  inv0d0 U1844 ( .I(n7661), .ZN(n3977) );
  inv0d0 U1846 ( .I(n6914), .ZN(n3941) );
  inv0d0 U1848 ( .I(n9428), .ZN(n3185) );
  inv0d0 U1850 ( .I(n5841), .ZN(n4746) );
  inv0d1 U1852 ( .I(n1355), .ZN(n1327) );
  inv0d1 U1854 ( .I(n1355), .ZN(n1328) );
  inv0d1 U1856 ( .I(n1123), .ZN(n1098) );
  inv0d1 U1857 ( .I(n1311), .ZN(n1276) );
  inv0d1 U1858 ( .I(n1312), .ZN(n1281) );
  inv0d1 U1859 ( .I(n1123), .ZN(n1099) );
  inv0d1 U1860 ( .I(n1355), .ZN(n1329) );
  inv0d1 U1924 ( .I(n1261), .ZN(n1234) );
  inv0d1 U1925 ( .I(n1312), .ZN(n1282) );
  inv0d1 U1958 ( .I(n1311), .ZN(n1277) );
  inv0d1 U1959 ( .I(n1312), .ZN(n1280) );
  inv0d1 U1960 ( .I(n1311), .ZN(n1274) );
  inv0d1 U1993 ( .I(n1355), .ZN(n1330) );
  inv0d0 U1994 ( .I(n8661), .ZN(n3219) );
  inv0d1 U1995 ( .I(n1260), .ZN(n1232) );
  inv0d1 U2028 ( .I(n1212), .ZN(n1189) );
  inv0d1 U2029 ( .I(n1165), .ZN(n1135) );
  inv0d1 U2030 ( .I(n1260), .ZN(n1228) );
  inv0d1 U2063 ( .I(n1212), .ZN(n1187) );
  inv0d1 U2064 ( .I(n1312), .ZN(n1279) );
  inv0d1 U2065 ( .I(n1261), .ZN(n1235) );
  inv0d1 U2098 ( .I(n1356), .ZN(n1326) );
  inv0d1 U2099 ( .I(n1312), .ZN(n1283) );
  inv0d1 U2100 ( .I(n1313), .ZN(n1289) );
  inv0d1 U2133 ( .I(n1166), .ZN(n1140) );
  inv0d1 U2134 ( .I(n1165), .ZN(n1138) );
  inv0d1 U2135 ( .I(n1122), .ZN(n1093) );
  inv0d1 U2136 ( .I(n1165), .ZN(n1136) );
  inv0d1 U2138 ( .I(n1165), .ZN(n1137) );
  inv0d1 U2139 ( .I(n1124), .ZN(n1100) );
  inv0d1 U2140 ( .I(n1123), .ZN(n1097) );
  inv0d1 U2174 ( .I(n1356), .ZN(n1325) );
  inv0d1 U2175 ( .I(n1124), .ZN(n1103) );
  inv0d1 U2273 ( .I(n1166), .ZN(n1141) );
  inv0d1 U2308 ( .I(n1124), .ZN(n1102) );
  inv0d1 U2309 ( .I(n1212), .ZN(n1190) );
  inv0d1 U2343 ( .I(n1260), .ZN(n1231) );
  inv0d1 U2378 ( .I(n1260), .ZN(n1229) );
  inv0d0 U2379 ( .I(n5773), .ZN(n3947) );
  inv0d1 U2381 ( .I(n1124), .ZN(n1104) );
  inv0d1 U2382 ( .I(n1311), .ZN(n1275) );
  inv0d0 U2384 ( .I(n8321), .ZN(n4019) );
  inv0d1 U2385 ( .I(n1166), .ZN(n1144) );
  inv0d1 U2387 ( .I(n1166), .ZN(n1139) );
  inv0d1 U2388 ( .I(n1311), .ZN(n1278) );
  inv0d1 U2390 ( .I(n1260), .ZN(n1233) );
  inv0d1 U2391 ( .I(n1166), .ZN(n1142) );
  inv0d1 U2393 ( .I(n1166), .ZN(n1143) );
  inv0d1 U2394 ( .I(n1125), .ZN(n1105) );
  inv0d1 U2396 ( .I(n1123), .ZN(n1094) );
  inv0d1 U2397 ( .I(n1212), .ZN(n1188) );
  inv0d0 U2399 ( .I(n10648), .ZN(n3942) );
  inv0d1 U2400 ( .I(n1313), .ZN(n1286) );
  inv0d1 U2402 ( .I(n1125), .ZN(n1106) );
  inv0d1 U2403 ( .I(n1261), .ZN(n1236) );
  inv0d1 U2405 ( .I(n1260), .ZN(n1230) );
  inv0d1 U2406 ( .I(n1313), .ZN(n1288) );
  inv0d1 U2408 ( .I(n1123), .ZN(n1096) );
  inv0d1 U2409 ( .I(n1123), .ZN(n1095) );
  inv0d1 U2411 ( .I(n1124), .ZN(n1101) );
  inv0d1 U2412 ( .I(n1313), .ZN(n1287) );
  inv0d0 U2414 ( .I(n7694), .ZN(n3887) );
  inv0d1 U2415 ( .I(n1355), .ZN(n1331) );
  inv0d1 U2417 ( .I(n1168), .ZN(n1149) );
  buffd1 U2418 ( .I(n696), .Z(n690) );
  buffd1 U2420 ( .I(n697), .Z(n689) );
  buffd1 U2421 ( .I(n697), .Z(n688) );
  buffd1 U2423 ( .I(n695), .Z(n694) );
  buffd1 U2424 ( .I(n695), .Z(n693) );
  buffd1 U2426 ( .I(n696), .Z(n692) );
  buffd1 U2427 ( .I(n696), .Z(n691) );
  buffd1 U2429 ( .I(n699), .Z(n682) );
  buffd1 U2430 ( .I(n700), .Z(n680) );
  buffd1 U2432 ( .I(n698), .Z(n686) );
  buffd1 U2433 ( .I(n698), .Z(n685) );
  buffd1 U2435 ( .I(n698), .Z(n684) );
  buffd1 U2436 ( .I(n699), .Z(n683) );
  buffd1 U2438 ( .I(n697), .Z(n687) );
  buffd1 U2439 ( .I(n699), .Z(n681) );
  buffd1 U2441 ( .I(n705), .Z(n665) );
  buffd1 U2442 ( .I(n704), .Z(n666) );
  buffd1 U2444 ( .I(n704), .Z(n668) );
  buffd1 U2445 ( .I(n704), .Z(n667) );
  buffd1 U2447 ( .I(n706), .Z(n660) );
  buffd1 U2448 ( .I(n706), .Z(n662) );
  buffd1 U2450 ( .I(n705), .Z(n663) );
  buffd1 U2451 ( .I(n705), .Z(n664) );
  buffd1 U2453 ( .I(n706), .Z(n661) );
  buffd1 U2454 ( .I(n701), .Z(n675) );
  buffd1 U2456 ( .I(n700), .Z(n678) );
  buffd1 U2457 ( .I(n701), .Z(n677) );
  buffd1 U2459 ( .I(n701), .Z(n676) );
  buffd1 U2460 ( .I(n703), .Z(n670) );
  buffd1 U2463 ( .I(n702), .Z(n672) );
  buffd1 U2464 ( .I(n702), .Z(n673) );
  buffd1 U2466 ( .I(n702), .Z(n674) );
  buffd1 U2467 ( .I(n703), .Z(n671) );
  buffd1 U2469 ( .I(n700), .Z(n679) );
  buffd1 U2470 ( .I(n703), .Z(n669) );
  inv0d0 U2472 ( .I(n8995), .ZN(n4190) );
  inv0d0 U2473 ( .I(n11762), .ZN(n3265) );
  inv0d1 U2475 ( .I(n1354), .ZN(n1332) );
  inv0d0 U2476 ( .I(n11626), .ZN(n3573) );
  inv0d1 U2478 ( .I(n1125), .ZN(n1110) );
  inv0d0 U2479 ( .I(n9565), .ZN(n2872) );
  inv0d0 U2481 ( .I(n7169), .ZN(n3278) );
  inv0d1 U2482 ( .I(n1168), .ZN(n1150) );
  inv0d1 U2484 ( .I(n1125), .ZN(n1107) );
  inv0d1 U2485 ( .I(n1312), .ZN(n1284) );
  inv0d1 U2486 ( .I(n1168), .ZN(n1151) );
  inv0d1 U2487 ( .I(n1125), .ZN(n1109) );
  inv0d1 U2488 ( .I(n1265), .ZN(n1256) );
  inv0d0 U2489 ( .I(n4774), .ZN(n3016) );
  inv0d1 U2490 ( .I(n1261), .ZN(n1237) );
  inv0d1 U2494 ( .I(n1313), .ZN(n1285) );
  inv0d1 U2495 ( .I(n1168), .ZN(n1152) );
  inv0d0 U2496 ( .I(n6320), .ZN(n3285) );
  inv0d1 U2498 ( .I(n1214), .ZN(n1194) );
  inv0d1 U2499 ( .I(n1125), .ZN(n1108) );
  inv0d1 U2501 ( .I(n1264), .ZN(n1250) );
  inv0d1 U2502 ( .I(n1216), .ZN(n1203) );
  inv0d1 U2503 ( .I(n1264), .ZN(n1251) );
  inv0d1 U2504 ( .I(n1317), .ZN(n1307) );
  inv0d1 U2505 ( .I(n1210), .ZN(n1178) );
  inv0d1 U2506 ( .I(n1127), .ZN(n1118) );
  inv0d1 U2507 ( .I(n1352), .ZN(n1348) );
  inv0d0 U2508 ( .I(n8637), .ZN(n3190) );
  inv0d1 U2509 ( .I(n1353), .ZN(n1343) );
  inv0d1 U2510 ( .I(n1210), .ZN(n1177) );
  inv0d1 U2511 ( .I(n1354), .ZN(n1333) );
  inv0d1 U2512 ( .I(n1261), .ZN(n1238) );
  inv0d1 U2513 ( .I(n1264), .ZN(n1252) );
  inv0d1 U2514 ( .I(n1216), .ZN(n1206) );
  inv0d1 U2515 ( .I(n1352), .ZN(n1347) );
  inv0d1 U2516 ( .I(n1352), .ZN(n1346) );
  inv0d1 U2517 ( .I(n1127), .ZN(n1119) );
  inv0d1 U2518 ( .I(n1264), .ZN(n1253) );
  inv0d1 U2519 ( .I(n1216), .ZN(n1204) );
  inv0d1 U2520 ( .I(n1354), .ZN(n1335) );
  inv0d1 U2521 ( .I(n1216), .ZN(n1205) );
  inv0d1 U2778 ( .I(n1168), .ZN(n1153) );
  inv0d1 U2780 ( .I(n1354), .ZN(n1334) );
  inv0d1 U2781 ( .I(n1317), .ZN(n1309) );
  inv0d1 U2783 ( .I(n1210), .ZN(n1179) );
  inv0d1 U2784 ( .I(n1265), .ZN(n1255) );
  inv0d1 U2785 ( .I(n1170), .ZN(n1163) );
  inv0d0 U2786 ( .I(n7370), .ZN(n3031) );
  inv0d1 U2788 ( .I(n1354), .ZN(n1336) );
  inv0d1 U2789 ( .I(n1170), .ZN(n1161) );
  inv0d1 U2793 ( .I(n1126), .ZN(n1111) );
  inv0d1 U2797 ( .I(n1317), .ZN(n1308) );
  inv0d1 U2799 ( .I(n1352), .ZN(n1345) );
  inv0d1 U2802 ( .I(n1352), .ZN(n1344) );
  inv0d1 U2804 ( .I(n1216), .ZN(n1207) );
  inv0d1 U2809 ( .I(n1265), .ZN(n1254) );
  inv0d0 U2828 ( .I(n11504), .ZN(n3993) );
  inv0d1 U2830 ( .I(n1354), .ZN(n1337) );
  inv0d1 U2832 ( .I(n1170), .ZN(n1162) );
  inv0d1 U2834 ( .I(n1167), .ZN(n1147) );
  inv0d1 U2842 ( .I(n1214), .ZN(n1195) );
  inv0d1 U2877 ( .I(n1353), .ZN(n1340) );
  inv0d1 U2883 ( .I(n1353), .ZN(n1339) );
  inv0d1 U2886 ( .I(n1126), .ZN(n1112) );
  inv0d1 U2889 ( .I(n1214), .ZN(n1198) );
  inv0d0 U2903 ( .I(n11985), .ZN(n3194) );
  inv0d1 U2911 ( .I(n1213), .ZN(n1191) );
  inv0d1 U2938 ( .I(n1214), .ZN(n1197) );
  inv0d1 U2944 ( .I(n1356), .ZN(n1324) );
  inv0d1 U2945 ( .I(n1168), .ZN(n1154) );
  inv0d1 U2946 ( .I(n1167), .ZN(n1146) );
  inv0d1 U2947 ( .I(n1214), .ZN(n1196) );
  inv0d1 U2952 ( .I(n1126), .ZN(n1116) );
  inv0d1 U2953 ( .I(n1122), .ZN(n1090) );
  inv0d1 U2954 ( .I(n1167), .ZN(n1145) );
  inv0d1 U2955 ( .I(n1127), .ZN(n1117) );
  inv0d1 U2957 ( .I(n1122), .ZN(n1092) );
  inv0d1 U2958 ( .I(n1126), .ZN(n1114) );
  inv0d1 U2960 ( .I(n1353), .ZN(n1341) );
  inv0d1 U2962 ( .I(n1353), .ZN(n1338) );
  inv0d1 U2963 ( .I(n1264), .ZN(n1249) );
  inv0d1 U2964 ( .I(n1212), .ZN(n1186) );
  inv0d1 U2965 ( .I(n1126), .ZN(n1113) );
  inv0d1 U2967 ( .I(n1213), .ZN(n1193) );
  inv0d1 U2968 ( .I(n1213), .ZN(n1192) );
  inv0d1 U2969 ( .I(n1122), .ZN(n1091) );
  inv0d0 U2970 ( .I(n5335), .ZN(n3708) );
  inv0d1 U2971 ( .I(n1126), .ZN(n1115) );
  inv0d0 U2973 ( .I(n6275), .ZN(n3389) );
  inv0d1 U2974 ( .I(n1167), .ZN(n1148) );
  inv0d0 U2975 ( .I(N5114), .ZN(n1396) );
  inv0d1 U2976 ( .I(n1353), .ZN(n1342) );
  inv0d0 U2977 ( .I(n9285), .ZN(n3428) );
  inv0d0 U2978 ( .I(n7774), .ZN(n3494) );
  inv0d0 U2979 ( .I(n6130), .ZN(n3523) );
  inv0d0 U2980 ( .I(n6803), .ZN(n4073) );
  inv0d0 U2981 ( .I(n6239), .ZN(n3358) );
  inv0d1 U2982 ( .I(n1314), .ZN(n1290) );
  inv0d0 U2983 ( .I(n9940), .ZN(n3738) );
  inv0d1 U2984 ( .I(n1164), .ZN(n1134) );
  inv0d1 U2985 ( .I(n1169), .ZN(n1155) );
  inv0d0 U2987 ( .I(n11402), .ZN(n4145) );
  inv0d0 U2988 ( .I(n5366), .ZN(n3543) );
  inv0d1 U2989 ( .I(n1314), .ZN(n1291) );
  inv0d0 U2990 ( .I(n9954), .ZN(n3769) );
  inv0d1 U2991 ( .I(n1315), .ZN(n1295) );
  inv0d0 U2992 ( .I(n5901), .ZN(n4123) );
  inv0d1 U2993 ( .I(n1215), .ZN(n1200) );
  inv0d1 U2994 ( .I(n1215), .ZN(n1199) );
  inv0d1 U2996 ( .I(n1351), .ZN(n1350) );
  inv0d1 U2997 ( .I(n1315), .ZN(n1298) );
  inv0d1 U2998 ( .I(n1169), .ZN(n1157) );
  inv0d1 U2999 ( .I(n1315), .ZN(n1296) );
  inv0d1 U3001 ( .I(n1351), .ZN(n1349) );
  inv0d1 U3002 ( .I(n1310), .ZN(n1272) );
  inv0d0 U3004 ( .I(n10369), .ZN(n2964) );
  inv0d1 U3007 ( .I(n1211), .ZN(n1184) );
  inv0d1 U3011 ( .I(n1316), .ZN(n1301) );
  inv0d1 U3012 ( .I(n1259), .ZN(n1226) );
  inv0d1 U3013 ( .I(n1211), .ZN(n1183) );
  inv0d1 U3015 ( .I(n1263), .ZN(n1248) );
  inv0d1 U3016 ( .I(n1211), .ZN(n1182) );
  inv0d1 U3017 ( .I(n1259), .ZN(n1225) );
  inv0d1 U3018 ( .I(n1315), .ZN(n1299) );
  inv0d1 U3020 ( .I(n1211), .ZN(n1181) );
  inv0d1 U3022 ( .I(n1316), .ZN(n1302) );
  inv0d1 U3023 ( .I(n1316), .ZN(n1303) );
  inv0d0 U3024 ( .I(n6522), .ZN(n2991) );
  inv0d1 U3026 ( .I(n1262), .ZN(n1242) );
  inv0d1 U3027 ( .I(n1169), .ZN(n1158) );
  inv0d1 U3037 ( .I(n1314), .ZN(n1293) );
  inv0d1 U3039 ( .I(n1263), .ZN(n1246) );
  inv0d1 U3046 ( .I(n1314), .ZN(n1292) );
  inv0d1 U3058 ( .I(n1121), .ZN(n1089) );
  inv0d1 U3079 ( .I(n1315), .ZN(n1297) );
  inv0d1 U3081 ( .I(n1316), .ZN(n1304) );
  inv0d1 U3091 ( .I(n1211), .ZN(n1180) );
  inv0d1 U3097 ( .I(n1215), .ZN(n1201) );
  inv0d0 U3105 ( .I(n6536), .ZN(n2972) );
  inv0d1 U3121 ( .I(n1316), .ZN(n1305) );
  inv0d1 U3138 ( .I(n1263), .ZN(n1247) );
  inv0d1 U3141 ( .I(n1263), .ZN(n1244) );
  inv0d1 U3145 ( .I(n1169), .ZN(n1159) );
  inv0d1 U3151 ( .I(n1314), .ZN(n1294) );
  inv0d1 U3156 ( .I(n1169), .ZN(n1156) );
  inv0d1 U3162 ( .I(n1262), .ZN(n1240) );
  inv0d1 U3168 ( .I(n1262), .ZN(n1239) );
  inv0d1 U3174 ( .I(n1262), .ZN(n1243) );
  inv0d1 U3180 ( .I(n1262), .ZN(n1241) );
  inv0d1 U3184 ( .I(n1263), .ZN(n1245) );
  inv0d0 U3188 ( .I(n10003), .ZN(n3549) );
  inv0d0 U3189 ( .I(n7114), .ZN(n3355) );
  inv0d0 U3197 ( .I(n4625), .ZN(n3252) );
  inv0d0 U3201 ( .I(n5149), .ZN(n3972) );
  inv0d0 U3206 ( .I(n11899), .ZN(n2836) );
  inv0d0 U3210 ( .I(n5677), .ZN(n2838) );
  inv0d0 U3214 ( .I(n11323), .ZN(n4587) );
  inv0d0 U3223 ( .I(n5039), .ZN(n4151) );
  inv0d0 U3226 ( .I(n6878), .ZN(n3917) );
  inv0d0 U3246 ( .I(n6361), .ZN(n3141) );
  inv0d0 U3247 ( .I(n8125), .ZN(n4374) );
  inv0d1 U3248 ( .I(n1217), .ZN(n1208) );
  inv0d0 U3249 ( .I(n8423), .ZN(n3857) );
  inv0d0 U3250 ( .I(n4861), .ZN(n2841) );
  inv0d0 U3251 ( .I(n7867), .ZN(n3267) );
  inv0d0 U3252 ( .I(n5975), .ZN(n4049) );
  inv0d0 U3253 ( .I(n4801), .ZN(n2933) );
  inv0d0 U3254 ( .I(n4431), .ZN(n3820) );
  inv0d0 U3256 ( .I(n11592), .ZN(n3672) );
  inv0d0 U3257 ( .I(n11601), .ZN(n3665) );
  inv0d1 U3260 ( .I(n1128), .ZN(n1120) );
  inv0d0 U3261 ( .I(n5317), .ZN(n3772) );
  inv0d0 U3262 ( .I(n9795), .ZN(n4077) );
  inv0d0 U3263 ( .I(n6644), .ZN(n4035) );
  inv0d0 U3266 ( .I(n6274), .ZN(n3357) );
  inv0d0 U3267 ( .I(n7178), .ZN(n3255) );
  inv0d0 U3268 ( .I(n6941), .ZN(n3824) );
  inv0d0 U3273 ( .I(n4707), .ZN(n3040) );
  inv0d0 U3274 ( .I(n10441), .ZN(n4766) );
  inv0d0 U3275 ( .I(n5015), .ZN(n4001) );
  inv0d0 U3276 ( .I(n7175), .ZN(n3280) );
  inv0d0 U3278 ( .I(n6951), .ZN(n3874) );
  inv0d0 U3279 ( .I(n7798), .ZN(n3499) );
  inv0d0 U3281 ( .I(n9602), .ZN(n3079) );
  inv0d0 U3284 ( .I(n7496), .ZN(n4232) );
  inv0d0 U3285 ( .I(n6632), .ZN(n3951) );
  inv0d0 U3286 ( .I(n7823), .ZN(n3403) );
  inv0d0 U3287 ( .I(n6047), .ZN(n3899) );
  inv0d0 U3291 ( .I(n8584), .ZN(n3260) );
  inv0d0 U3292 ( .I(N13650), .ZN(n7604) );
  inv0d0 U3293 ( .I(n1724), .ZN(N13650) );
  inv0d0 U3294 ( .I(n6129), .ZN(n3520) );
  inv0d0 U3295 ( .I(n5965), .ZN(n4012) );
  inv0d0 U3298 ( .I(n10271), .ZN(n2975) );
  inv0d0 U3299 ( .I(n7256), .ZN(n3145) );
  inv0d0 U3300 ( .I(n988), .ZN(n983) );
  inv0d0 U3302 ( .I(N3182), .ZN(n419) );
  oaim21d1 U3303 ( .B1(n2754), .B2(n3589), .A(n2753), .ZN(n3594) );
  nr02d1 U3306 ( .A1(n2777), .A2(n3617), .ZN(n3622) );
  inv0d0 U3309 ( .I(n3655), .ZN(n2770) );
  oaim21d1 U3312 ( .B1(n3648), .B2(n3589), .A(n2753), .ZN(n3623) );
  nr02d1 U3315 ( .A1(n503), .A2(N3179), .ZN(n402) );
  inv0d0 U3317 ( .I(n496), .ZN(n2756) );
  nr02d1 U3318 ( .A1(n505), .A2(N3976), .ZN(n385) );
  an02d1 U3319 ( .A1(n3649), .A2(n3647), .Z(n3583) );
  nr02d1 U3320 ( .A1(N3976), .A2(N3179), .ZN(n404) );
  inv0d0 U3321 ( .I(n2709), .ZN(n2721) );
  inv0d0 U3322 ( .I(n3651), .ZN(n2775) );
  inv0d0 U3323 ( .I(n3707), .ZN(n2758) );
  buffd1 U3324 ( .I(n3797), .Z(n937) );
  buffd1 U3325 ( .I(n3797), .Z(n938) );
  buffd1 U3327 ( .I(n3797), .Z(n939) );
  buffd1 U3328 ( .I(n3797), .Z(n940) );
  buffd1 U3329 ( .I(n3710), .Z(n945) );
  buffd1 U3330 ( .I(n3710), .Z(n947) );
  buffd1 U3331 ( .I(n3710), .Z(n946) );
  buffd1 U3334 ( .I(n4131), .Z(n893) );
  buffd1 U3336 ( .I(n4100), .Z(n897) );
  buffd1 U3339 ( .I(n4069), .Z(n901) );
  buffd1 U3340 ( .I(n4040), .Z(n905) );
  buffd1 U3341 ( .I(n4162), .Z(n890) );
  buffd1 U3344 ( .I(n4131), .Z(n894) );
  buffd1 U3345 ( .I(n4100), .Z(n898) );
  buffd1 U3347 ( .I(n3980), .Z(n914) );
  buffd1 U3348 ( .I(n4194), .Z(n886) );
  buffd1 U3350 ( .I(n3980), .Z(n915) );
  buffd1 U3351 ( .I(n4194), .Z(n885) );
  buffd1 U3352 ( .I(n4162), .Z(n889) );
  buffd1 U3353 ( .I(n4069), .Z(n902) );
  buffd1 U3354 ( .I(n4131), .Z(n895) );
  buffd1 U3355 ( .I(n4011), .Z(n911) );
  buffd1 U3357 ( .I(n3980), .Z(n913) );
  buffd1 U3358 ( .I(n4100), .Z(n899) );
  buffd1 U3359 ( .I(n4069), .Z(n903) );
  buffd1 U3361 ( .I(n4040), .Z(n907) );
  buffd1 U3362 ( .I(n4040), .Z(n906) );
  buffd1 U3366 ( .I(n4011), .Z(n910) );
  buffd1 U3382 ( .I(n4194), .Z(n887) );
  buffd1 U3386 ( .I(n4011), .Z(n909) );
  buffd1 U3391 ( .I(n4162), .Z(n891) );
  buffd1 U3408 ( .I(n3710), .Z(n948) );
  buffd1 U3415 ( .I(n4162), .Z(n892) );
  buffd1 U3419 ( .I(n4100), .Z(n900) );
  buffd1 U3424 ( .I(n4069), .Z(n904) );
  buffd1 U3426 ( .I(n4011), .Z(n912) );
  buffd1 U3427 ( .I(n3980), .Z(n916) );
  buffd1 U3439 ( .I(n4131), .Z(n896) );
  buffd1 U3446 ( .I(n4040), .Z(n908) );
  buffd1 U3449 ( .I(n4194), .Z(n888) );
  buffd1 U3453 ( .I(n3949), .Z(n917) );
  buffd1 U3455 ( .I(n3885), .Z(n925) );
  buffd1 U3461 ( .I(n3949), .Z(n918) );
  buffd1 U3463 ( .I(n3918), .Z(n922) );
  buffd1 U3470 ( .I(n3885), .Z(n926) );
  buffd1 U3472 ( .I(n3949), .Z(n919) );
  buffd1 U3481 ( .I(n3855), .Z(n931) );
  buffd1 U3489 ( .I(n3827), .Z(n935) );
  buffd1 U3492 ( .I(n3855), .Z(n929) );
  buffd1 U3498 ( .I(n3827), .Z(n933) );
  buffd1 U3511 ( .I(n3767), .Z(n941) );
  buffd1 U3514 ( .I(n3918), .Z(n923) );
  buffd1 U3527 ( .I(n3918), .Z(n921) );
  buffd1 U3528 ( .I(n3767), .Z(n942) );
  buffd1 U3535 ( .I(n3885), .Z(n927) );
  buffd1 U3542 ( .I(n3767), .Z(n943) );
  buffd1 U3545 ( .I(n3855), .Z(n930) );
  buffd1 U3546 ( .I(n3827), .Z(n934) );
  inv0d0 U3548 ( .I(n3662), .ZN(n2766) );
  buffd1 U3560 ( .I(n3918), .Z(n924) );
  buffd1 U3569 ( .I(n3885), .Z(n928) );
  buffd1 U3571 ( .I(n3855), .Z(n932) );
  buffd1 U3583 ( .I(n3827), .Z(n936) );
  buffd1 U3598 ( .I(n3949), .Z(n920) );
  buffd1 U3607 ( .I(n3767), .Z(n944) );
  nd02d1 U3611 ( .A1(n2771), .A2(n493), .ZN(n3667) );
  buffd1 U3613 ( .I(n738), .Z(n740) );
  buffd1 U3618 ( .I(n738), .Z(n741) );
  buffd1 U3623 ( .I(n738), .Z(n742) );
  buffd1 U3630 ( .I(n754), .Z(n756) );
  buffd1 U3633 ( .I(n754), .Z(n757) );
  buffd1 U3635 ( .I(n754), .Z(n758) );
  inv0d0 U3639 ( .I(n2), .ZN(n2768) );
  buffd1 U3641 ( .I(n773), .Z(n775) );
  buffd1 U3642 ( .I(n773), .Z(n776) );
  buffd1 U3643 ( .I(n773), .Z(n777) );
  buffd1 U3644 ( .I(n797), .Z(n799) );
  buffd1 U3645 ( .I(n797), .Z(n800) );
  buffd1 U3646 ( .I(n797), .Z(n801) );
  buffd1 U3647 ( .I(n767), .Z(n769) );
  buffd1 U3648 ( .I(n767), .Z(n770) );
  buffd1 U3651 ( .I(n767), .Z(n771) );
  buffd1 U3655 ( .I(n712), .Z(n714) );
  buffd1 U3659 ( .I(n712), .Z(n715) );
  buffd1 U3661 ( .I(n712), .Z(n716) );
  buffd1 U3662 ( .I(n725), .Z(n727) );
  buffd1 U3666 ( .I(n725), .Z(n728) );
  buffd1 U3669 ( .I(n725), .Z(n729) );
  buffd1 U3677 ( .I(n810), .Z(n812) );
  buffd1 U3678 ( .I(n810), .Z(n813) );
  buffd1 U3680 ( .I(n810), .Z(n814) );
  inv0d0 U3681 ( .I(N3181), .ZN(n418) );
  buffd1 U3682 ( .I(n4335), .Z(n838) );
  buffd1 U3683 ( .I(n4335), .Z(n839) );
  nd02d1 U3684 ( .A1(n4345), .A2(n495), .ZN(n4343) );
  buffd1 U3687 ( .I(n4327), .Z(n857) );
  buffd1 U3689 ( .I(n4327), .Z(n856) );
  buffd1 U3690 ( .I(n4327), .Z(n855) );
  nd02d1 U3691 ( .A1(n495), .A2(n2781), .ZN(n4258) );
  buffd1 U3692 ( .I(n4327), .Z(n858) );
  buffd1 U3693 ( .I(n4364), .Z(n744) );
  buffd1 U3694 ( .I(n4364), .Z(n745) );
  nd02d1 U3696 ( .A1(n4345), .A2(n2), .ZN(n4371) );
  nd02d1 U3698 ( .A1(n2), .A2(n2781), .ZN(n4354) );
  buffd1 U3699 ( .I(n4327), .Z(n860) );
  buffd1 U3700 ( .I(n4327), .Z(n859) );
  buffd1 U3702 ( .I(n4327), .Z(n861) );
  buffd1 U3704 ( .I(n840), .Z(n847) );
  buffd1 U3710 ( .I(n4335), .Z(n840) );
  buffd1 U3711 ( .I(n4358), .Z(n779) );
  buffd1 U3712 ( .I(n4358), .Z(n780) );
  buffd1 U3716 ( .I(n4358), .Z(n781) );
  buffd1 U3717 ( .I(n746), .Z(n753) );
  buffd1 U3718 ( .I(n4364), .Z(n746) );
  buffd1 U3719 ( .I(n3671), .Z(n497) );
  nr02d1 U3721 ( .A1(n3667), .A2(n2777), .ZN(n3671) );
  nd02d1 U3722 ( .A1(n3647), .A2(n2771), .ZN(n3590) );
  inv0d0 U3724 ( .I(n1384), .ZN(n1403) );
  inv0d0 U3725 ( .I(n1390), .ZN(n1401) );
  inv0d0 U3726 ( .I(n1381), .ZN(n1402) );
  nd03d1 U3727 ( .A1(n4949), .A2(n5837), .A3(n5427), .ZN(n12048) );
  nr02d1 U3729 ( .A1(n7333), .A2(n4839), .ZN(n7987) );
  nr02d1 U3730 ( .A1(n3382), .A2(n6252), .ZN(n7135) );
  nd02d1 U3731 ( .A1(n10329), .A2(n2889), .ZN(n4904) );
  inv0d0 U3732 ( .I(n2527), .ZN(N8840) );
  inv0d0 U3733 ( .I(n5545), .ZN(n3209) );
  inv0d0 U3734 ( .I(n11766), .ZN(n3307) );
  inv0d0 U3735 ( .I(n4943), .ZN(n3096) );
  inv0d0 U3736 ( .I(n1477), .ZN(n1479) );
  nd02d1 U3737 ( .A1(N14562), .A2(n8730), .ZN(n6557) );
  nd03d1 U3739 ( .A1(n5042), .A2(n4196), .A3(n4078), .ZN(n5038) );
  nd02d1 U3740 ( .A1(n4391), .A2(n3932), .ZN(n4387) );
  nr02d1 U3742 ( .A1(n8836), .A2(n3206), .ZN(n11806) );
  inv0d0 U3744 ( .I(n2002), .ZN(N11858) );
  inv0d0 U3745 ( .I(n5736), .ZN(n3512) );
  inv0d0 U3747 ( .I(n5371), .ZN(n3550) );
  nd02d1 U3750 ( .A1(N14178), .A2(n3050), .ZN(n6577) );
  nd02d1 U3751 ( .A1(N10461), .A2(n9139), .ZN(n7428) );
  nd03d1 U3752 ( .A1(n5093), .A2(n5777), .A3(n11536), .ZN(n11541) );
  nr02d1 U3754 ( .A1(n4601), .A2(n7381), .ZN(n6314) );
  inv0d0 U3758 ( .I(n11815), .ZN(n3147) );
  inv0d0 U3763 ( .I(n4932), .ZN(n2832) );
  inv0d0 U3767 ( .I(n9370), .ZN(n3261) );
  nr02d1 U3768 ( .A1(n6281), .A2(n6275), .ZN(n8581) );
  nd02d1 U3771 ( .A1(n3999), .A2(n4000), .ZN(n5041) );
  aoim22d1 U3775 ( .A1(n3071), .A2(n5596), .B1(n5597), .B2(n5598), .Z(n5594)
         );
  nr02d1 U3776 ( .A1(n9315), .A2(n11242), .ZN(n5416) );
  inv0d0 U3777 ( .I(n8061), .ZN(n3176) );
  inv0d0 U3778 ( .I(n4630), .ZN(n3304) );
  nd02d1 U3779 ( .A1(n3265), .A2(n4627), .ZN(n11768) );
  nr02d1 U3782 ( .A1(n6584), .A2(n7258), .ZN(n9453) );
  nd12d1 U3784 ( .A1(n1730), .A2(n11779), .ZN(n6365) );
  nd03d1 U3786 ( .A1(n8802), .A2(n2861), .A3(n8798), .ZN(n4863) );
  nr02d1 U3787 ( .A1(n7011), .A2(n5339), .ZN(n6111) );
  nr02d1 U3788 ( .A1(n9935), .A2(n6059), .ZN(n6062) );
  inv0d0 U3789 ( .I(n1985), .ZN(n1988) );
  nd02d1 U3794 ( .A1(N11256), .A2(n11605), .ZN(n6987) );
  nd02d1 U3803 ( .A1(N11618), .A2(n10402), .ZN(n8464) );
  nd02d1 U3824 ( .A1(n11208), .A2(n3010), .ZN(n8744) );
  nd12d1 U3831 ( .A1(n1889), .A2(n3362), .ZN(n6198) );
  nr02d1 U3835 ( .A1(n7385), .A2(n7169), .ZN(n5480) );
  nd02d1 U3839 ( .A1(N13858), .A2(n7227), .ZN(n7236) );
  inv0d0 U3844 ( .I(n1698), .ZN(N13858) );
  inv0d0 U3855 ( .I(n1697), .ZN(n1699) );
  nr02d1 U3861 ( .A1(n10285), .A2(n10282), .ZN(n11126) );
  nd02d1 U3864 ( .A1(N15186), .A2(n8831), .ZN(n7337) );
  nd02d1 U3868 ( .A1(N14210), .A2(n6442), .ZN(n6448) );
  nd03d1 U3875 ( .A1(n4034), .A2(n8340), .A3(n10617), .ZN(n10414) );
  nd02d1 U3878 ( .A1(n3446), .A2(n3421), .ZN(n6188) );
  nd02d1 U3883 ( .A1(N10041), .A2(n8340), .ZN(n8337) );
  nd02d1 U3887 ( .A1(N14194), .A2(n10172), .ZN(n8688) );
  inv0d0 U3888 ( .I(n1644), .ZN(n1647) );
  nr02d1 U3894 ( .A1(n6353), .A2(n6347), .ZN(n8839) );
  nr02d1 U3896 ( .A1(n4995), .A2(n8520), .ZN(n8528) );
  nd02d1 U3904 ( .A1(n8340), .A2(n9846), .ZN(n8344) );
  inv0d0 U3907 ( .I(n5525), .ZN(n3181) );
  nd03d1 U3912 ( .A1(n8857), .A2(n7003), .A3(n5544), .ZN(n5750) );
  nd02d1 U3915 ( .A1(N14066), .A2(n8670), .ZN(n11009) );
  nd02d1 U3917 ( .A1(n9601), .A2(n3115), .ZN(n6564) );
  nr02d1 U3919 ( .A1(n6690), .A2(n6686), .ZN(n5796) );
  nd03d1 U3921 ( .A1(n3013), .A2(n11854), .A3(N14626), .ZN(n7973) );
  nd02d1 U3924 ( .A1(n4960), .A2(n3234), .ZN(n5552) );
  nd02d1 U3932 ( .A1(N14482), .A2(n11978), .ZN(n6478) );
  nd02d1 U3934 ( .A1(n2950), .A2(n8047), .ZN(n7313) );
  nd02d1 U3938 ( .A1(n3841), .A2(n10683), .ZN(n4409) );
  nd02d1 U3942 ( .A1(N13906), .A2(n11983), .ZN(n9437) );
  nd02d1 U3944 ( .A1(N13266), .A2(n7384), .ZN(n7169) );
  inv0d0 U3956 ( .I(n1777), .ZN(n1780) );
  nd02d1 U3964 ( .A1(n9104), .A2(n5077), .ZN(n6860) );
  nd02d1 U3967 ( .A1(n12059), .A2(n5767), .ZN(n6016) );
  nd03d1 U3974 ( .A1(n5314), .A2(n5794), .A3(n9651), .ZN(n7461) );
  nd02d1 U3977 ( .A1(N13058), .A2(n5463), .ZN(n6275) );
  oai311d1 U3982 ( .C1(n1229), .C2(n1178), .C3(n1701), .A(n1297), .B(n1335), 
        .ZN(n14) );
  nd02d1 U3983 ( .A1(n9502), .A2(n3008), .ZN(n8030) );
  nd02d1 U3989 ( .A1(N9554), .A2(n4093), .ZN(n6830) );
  nd03d1 U3992 ( .A1(n6079), .A2(n2849), .A3(N15170), .ZN(n7335) );
  nd02d1 U3999 ( .A1(N15090), .A2(n8783), .ZN(n10357) );
  nd02d1 U4000 ( .A1(N13586), .A2(n3169), .ZN(n7211) );
  nd02d1 U4002 ( .A1(N14802), .A2(n2957), .ZN(n7315) );
  nd02d1 U4006 ( .A1(N13298), .A2(n11752), .ZN(n4601) );
  nd02d1 U4008 ( .A1(N12546), .A2(n9319), .ZN(n5418) );
  nd02d1 U4016 ( .A1(n11779), .A2(n3166), .ZN(n5510) );
  nd02d1 U4021 ( .A1(n3125), .A2(n7939), .ZN(n6459) );
  nd02d1 U4033 ( .A1(N12594), .A2(n12018), .ZN(n6197) );
  inv0d0 U4034 ( .I(n1888), .ZN(N12594) );
  nd02d1 U4042 ( .A1(N14418), .A2(n3116), .ZN(n7963) );
  nd03d1 U4046 ( .A1(n4972), .A2(n5044), .A3(n7187), .ZN(n7201) );
  nd02d1 U4058 ( .A1(n11779), .A2(n3167), .ZN(n7214) );
  nd02d1 U4059 ( .A1(n11830), .A2(n3127), .ZN(n5583) );
  nr02d1 U4062 ( .A1(n4713), .A2(n3050), .ZN(n4710) );
  nd02d1 U4063 ( .A1(N15538), .A2(n10329), .ZN(n11954) );
  nd02d1 U4067 ( .A1(n4945), .A2(n3115), .ZN(n11053) );
  nd03d1 U4069 ( .A1(n5140), .A2(n4950), .A3(n7276), .ZN(n7281) );
  nd12d1 U4071 ( .A1(n1749), .A2(n6333), .ZN(n5500) );
  nr02d1 U4072 ( .A1(n10307), .A2(n10297), .ZN(n11137) );
  nd02d1 U4075 ( .A1(n3943), .A2(n9139), .ZN(n4433) );
  nd03d1 U4076 ( .A1(n6665), .A2(n5778), .A3(n6666), .ZN(n5820) );
  nd02d1 U4077 ( .A1(N15378), .A2(n2882), .ZN(n11186) );
  nd02d1 U4078 ( .A1(N14498), .A2(n3112), .ZN(n6487) );
  nd02d1 U4082 ( .A1(N13682), .A2(n10969), .ZN(n8620) );
  nd02d1 U4083 ( .A1(n5652), .A2(n3807), .ZN(n10722) );
  nd02d1 U4087 ( .A1(n2914), .A2(n11898), .ZN(n10280) );
  nd02d1 U4088 ( .A1(n2831), .A2(n10359), .ZN(n4850) );
  inv0d0 U4089 ( .I(n4722), .ZN(n3022) );
  nd02d1 U4091 ( .A1(n3035), .A2(n6430), .ZN(n7370) );
  nd02d1 U4094 ( .A1(N11151), .A2(n6976), .ZN(n5286) );
  inv0d0 U4095 ( .I(n2097), .ZN(n2099) );
  nr02d1 U4097 ( .A1(n8801), .A2(n8798), .ZN(n11962) );
  nd02d1 U4098 ( .A1(N8025), .A2(n11304), .ZN(n9652) );
  nd02d1 U4100 ( .A1(n3110), .A2(n3111), .ZN(n6480) );
  nd02d1 U4102 ( .A1(N14578), .A2(n3104), .ZN(n4778) );
  nd02d1 U4104 ( .A1(N13346), .A2(n3289), .ZN(n10097) );
  nd02d1 U4107 ( .A1(N11061), .A2(n3810), .ZN(n6059) );
  nd02d1 U4108 ( .A1(n11893), .A2(n2914), .ZN(n4932) );
  nd03d1 U4110 ( .A1(n5751), .A2(n5182), .A3(n6983), .ZN(n6996) );
  nr02d1 U4112 ( .A1(n9071), .A2(n5940), .ZN(n6821) );
  nd12d1 U4113 ( .A1(n1789), .A2(n4592), .ZN(n7857) );
  nd03d1 U4114 ( .A1(n3471), .A2(n3469), .A3(n3470), .ZN(n4495) );
  nr02d1 U4115 ( .A1(n8620), .A2(n8621), .ZN(n7216) );
  nd02d1 U4120 ( .A1(n6746), .A2(n6666), .ZN(n6741) );
  nd03d1 U4121 ( .A1(n11333), .A2(n7487), .A3(N8282), .ZN(n9687) );
  nd02d1 U4123 ( .A1(N12162), .A2(n5384), .ZN(n5388) );
  nd02d1 U4124 ( .A1(n11840), .A2(n3120), .ZN(n10382) );
  nd02d1 U4125 ( .A1(n11304), .A2(n8897), .ZN(n8893) );
  nd02d1 U4126 ( .A1(n11220), .A2(n3204), .ZN(n7898) );
  nd02d1 U4128 ( .A1(N14242), .A2(n3126), .ZN(n7948) );
  nd02d1 U4129 ( .A1(N13410), .A2(n10099), .ZN(n4623) );
  nr02d1 U4131 ( .A1(n8190), .A2(n7458), .ZN(n5788) );
  nd02d1 U4132 ( .A1(N11730), .A2(n9977), .ZN(n7031) );
  nd02d1 U4133 ( .A1(n7605), .A2(n3991), .ZN(n7610) );
  aoim22d1 U4134 ( .A1(n7697), .A2(n11576), .B1(n6043), .B2(n11577), .Z(n11575) );
  nr02d1 U4135 ( .A1(n6165), .A2(n9268), .ZN(n5368) );
  nr02d1 U4139 ( .A1(n5999), .A2(n9139), .ZN(n5172) );
  nd02d1 U4140 ( .A1(N10686), .A2(n5201), .ZN(n6029) );
  nr02d1 U4143 ( .A1(n11755), .A2(n5520), .ZN(n11757) );
  nd02d1 U4144 ( .A1(n4392), .A2(n5870), .ZN(n11330) );
  nd02d1 U4145 ( .A1(n8524), .A2(n4439), .ZN(n4995) );
  nd03d1 U4146 ( .A1(n4006), .A2(n4056), .A3(N9696), .ZN(n5050) );
  nd02d1 U4147 ( .A1(n11208), .A2(n11850), .ZN(n4788) );
  nr02d1 U4149 ( .A1(n5500), .A2(n5501), .ZN(n10953) );
  nd02d1 U4150 ( .A1(n4039), .A2(n6640), .ZN(n8343) );
  nd03d1 U4152 ( .A1(n5795), .A2(n5796), .A3(n4261), .ZN(n5792) );
  inv0d0 U4154 ( .I(n5310), .ZN(n3771) );
  nd02d1 U4155 ( .A1(n6351), .A2(n3146), .ZN(n6361) );
  nr02d1 U4158 ( .A1(n5475), .A2(n5474), .ZN(n7850) );
  nd03d1 U4160 ( .A1(n10825), .A2(n12022), .A3(n3431), .ZN(n4502) );
  nd02d1 U4161 ( .A1(n2932), .A2(n4938), .ZN(n4831) );
  nd02d1 U4162 ( .A1(N9456), .A2(n4083), .ZN(n5017) );
  nd02d1 U4164 ( .A1(n6936), .A2(n3956), .ZN(n5187) );
  nd12d1 U4165 ( .A1(n15), .A2(n7311), .ZN(n8756) );
  nd04d1 U4172 ( .A1(n1341), .A2(n1299), .A3(n1247), .A4(n1546), .ZN(n15) );
  nd03d1 U4174 ( .A1(n5895), .A2(n4116), .A3(n5886), .ZN(n5019) );
  inv0d0 U4176 ( .I(n4678), .ZN(n3203) );
  inv0d0 U4178 ( .I(n5559), .ZN(n3212) );
  nd02d1 U4182 ( .A1(n3272), .A2(n8581), .ZN(n4579) );
  nd02d1 U4184 ( .A1(N10761), .A2(n3845), .ZN(n5214) );
  nr02d1 U4186 ( .A1(n4920), .A2(n11937), .ZN(n4888) );
  nd12d1 U4187 ( .A1(n16), .A2(n2967), .ZN(n10366) );
  nd04d1 U4188 ( .A1(n1342), .A2(n1300), .A3(n1247), .A4(n1531), .ZN(n16) );
  nd02d1 U4190 ( .A1(n3103), .A2(n3104), .ZN(n8726) );
  nd02d1 U4191 ( .A1(N9624), .A2(n4057), .ZN(n5951) );
  nd02d1 U4197 ( .A1(N14162), .A2(n8680), .ZN(n10386) );
  nd02d1 U4198 ( .A1(n3112), .A2(n3090), .ZN(n4763) );
  nd02d1 U4199 ( .A1(N9846), .A2(n9104), .ZN(n9100) );
  nd02d1 U4200 ( .A1(N15026), .A2(n11968), .ZN(n4840) );
  nd02d1 U4203 ( .A1(n7356), .A2(n2979), .ZN(n6542) );
  nr02d1 U4205 ( .A1(n10393), .A2(n11708), .ZN(n4548) );
  nd02d1 U4206 ( .A1(n6936), .A2(n3828), .ZN(n4431) );
  nd02d1 U4207 ( .A1(n8193), .A2(n6719), .ZN(n8203) );
  nr02d1 U4208 ( .A1(n8626), .A2(n10126), .ZN(n11791) );
  nd02d1 U4210 ( .A1(N13986), .A2(n3234), .ZN(n6406) );
  nd03d1 U4213 ( .A1(n4262), .A2(n4266), .A3(n4268), .ZN(n6730) );
  nd03d1 U4219 ( .A1(n5271), .A2(n5433), .A3(n8414), .ZN(n8430) );
  nd03d1 U4220 ( .A1(n4949), .A2(n5427), .A3(n6114), .ZN(n6118) );
  inv0d0 U4221 ( .I(n5657), .ZN(n2963) );
  nr02d1 U4222 ( .A1(n7963), .A2(n11839), .ZN(n7362) );
  nd02d1 U4223 ( .A1(N14258), .A2(n3061), .ZN(n7935) );
  nd02d1 U4224 ( .A1(n10882), .A2(n6232), .ZN(n6237) );
  nd02d1 U4225 ( .A1(n11208), .A2(n8030), .ZN(n11850) );
  nr02d1 U4226 ( .A1(n9718), .A2(n8215), .ZN(n6727) );
  nd02d1 U4227 ( .A1(n7206), .A2(n3146), .ZN(n7210) );
  nd02d1 U4228 ( .A1(N13538), .A2(n8838), .ZN(n6347) );
  nd02d1 U4229 ( .A1(n11968), .A2(n9539), .ZN(n11966) );
  nd03d1 U4230 ( .A1(n5904), .A2(n11833), .A3(N14402), .ZN(n11047) );
  nd03d1 U4231 ( .A1(n5621), .A2(n8691), .A3(N14306), .ZN(n6460) );
  nr02d1 U4233 ( .A1(n9981), .A2(n7031), .ZN(n5744) );
  nd03d1 U4236 ( .A1(N9092), .A2(n4169), .A3(N9106), .ZN(n9769) );
  inv0d0 U4237 ( .I(n7881), .ZN(n3153) );
  inv0d0 U4251 ( .I(n7886), .ZN(n3154) );
  nd02d1 U4255 ( .A1(n4296), .A2(n4281), .ZN(n6671) );
  nd02d1 U4257 ( .A1(N14946), .A2(n11970), .ZN(n10258) );
  nd02d1 U4259 ( .A1(N14098), .A2(n6430), .ZN(n6440) );
  nr02d1 U4283 ( .A1(n7211), .A2(n3167), .ZN(n9607) );
  nd02d1 U4286 ( .A1(n3545), .A2(n9255), .ZN(n9261) );
  nd02d1 U4290 ( .A1(N11496), .A2(n8453), .ZN(n5339) );
  nd03d1 U4293 ( .A1(n7423), .A2(n5181), .A3(n3977), .ZN(n8086) );
  nr02d1 U4301 ( .A1(n7760), .A2(n4449), .ZN(n7759) );
  nd02d1 U4308 ( .A1(N11376), .A2(n11615), .ZN(n5319) );
  nd02d1 U4313 ( .A1(n4441), .A2(n5001), .ZN(n4467) );
  inv0d0 U4336 ( .I(n9651), .ZN(n2773) );
  inv0d0 U4340 ( .I(n9653), .ZN(n2810) );
  nd03d1 U4345 ( .A1(n9081), .A2(n4966), .A3(N9610), .ZN(n6834) );
  nd02d1 U4349 ( .A1(n3509), .A2(n5001), .ZN(n11649) );
  nd02d1 U4352 ( .A1(n5865), .A2(n6660), .ZN(n5871) );
  nd02d1 U4355 ( .A1(N13730), .A2(n8624), .ZN(n6377) );
  nd03d1 U4356 ( .A1(n4376), .A2(n11336), .A3(n4384), .ZN(n8125) );
  nd02d1 U4359 ( .A1(N9652), .A2(n4003), .ZN(n5015) );
  nd02d1 U4368 ( .A1(N14738), .A2(n3006), .ZN(n9512) );
  nd03d1 U4382 ( .A1(n4106), .A2(n12065), .A3(N9442), .ZN(n7581) );
  nd02d1 U4388 ( .A1(N14370), .A2(n11833), .ZN(n10188) );
  nd02d1 U4394 ( .A1(n9624), .A2(n3774), .ZN(n5317) );
  nd02d1 U4399 ( .A1(N13506), .A2(n5718), .ZN(n5512) );
  nd02d1 U4407 ( .A1(N12514), .A2(n3445), .ZN(n10847) );
  nd03d1 U4409 ( .A1(n4086), .A2(n4102), .A3(N9484), .ZN(n7590) );
  nd02d1 U4414 ( .A1(N12914), .A2(n6247), .ZN(n6254) );
  nd02d1 U4416 ( .A1(n2909), .A2(n2879), .ZN(n8821) );
  nd02d1 U4417 ( .A1(N15410), .A2(n11931), .ZN(n10350) );
  nd02d1 U4421 ( .A1(n2966), .A2(n2964), .ZN(n7357) );
  nd02d1 U4426 ( .A1(n3293), .A2(n7189), .ZN(n5492) );
  nd02d1 U4427 ( .A1(N13234), .A2(n10918), .ZN(n7386) );
  nd03d1 U4433 ( .A1(n4961), .A2(n4960), .A3(n3140), .ZN(n5551) );
  nd02d1 U4435 ( .A1(n7227), .A2(n3189), .ZN(n4667) );
  nr02d1 U4443 ( .A1(n11568), .A2(n5216), .ZN(n11572) );
  inv0d0 U4447 ( .I(n4898), .ZN(n2891) );
  nd02d1 U4454 ( .A1(N14594), .A2(n11854), .ZN(n8731) );
  nd03d1 U4455 ( .A1(n5852), .A2(n6661), .A3(n5847), .ZN(n5856) );
  nd02d1 U4457 ( .A1(n3041), .A2(n3050), .ZN(n4707) );
  nd03d1 U4469 ( .A1(n5101), .A2(n5082), .A3(n5085), .ZN(n5089) );
  nd03d1 U4470 ( .A1(n4271), .A2(n6719), .A3(N8549), .ZN(n9714) );
  nd02d1 U4473 ( .A1(N10161), .A2(n3967), .ZN(n5123) );
  nd02d1 U4477 ( .A1(n4897), .A2(n4917), .ZN(n4896) );
  inv0d0 U4483 ( .I(n9333), .ZN(n3410) );
  inv0d0 U4491 ( .I(n6226), .ZN(n3409) );
  nd02d1 U4494 ( .A1(n3060), .A2(n3061), .ZN(n9468) );
  nd02d1 U4496 ( .A1(N9666), .A2(n11473), .ZN(n5006) );
  nd02d1 U4497 ( .A1(n8838), .A2(n3300), .ZN(n8616) );
  nd02d1 U4501 ( .A1(N11391), .A2(n3778), .ZN(n10734) );
  nd02d1 U4502 ( .A1(n6521), .A2(n4938), .ZN(n6534) );
  nd02d1 U4507 ( .A1(n4826), .A2(n10257), .ZN(n4837) );
  nd02d1 U4508 ( .A1(N11466), .A2(n3787), .ZN(n5334) );
  nd02d1 U4509 ( .A1(n5567), .A2(n9879), .ZN(n6914) );
  nd02d1 U4510 ( .A1(N15458), .A2(n11937), .ZN(n11155) );
  nd02d1 U4511 ( .A1(n5567), .A2(n5096), .ZN(n6634) );
  nd02d1 U4512 ( .A1(n5163), .A2(n3936), .ZN(n5158) );
  nd02d1 U4513 ( .A1(N11091), .A2(n3736), .ZN(n6066) );
  nd02d1 U4514 ( .A1(N11121), .A2(n8433), .ZN(n5279) );
  nd02d1 U4516 ( .A1(n4092), .A2(n8876), .ZN(n6829) );
  nd02d1 U4518 ( .A1(n4115), .A2(n5293), .ZN(n6786) );
  nd02d1 U4519 ( .A1(n5245), .A2(n5758), .ZN(n5251) );
  nd02d1 U4521 ( .A1(n7472), .A2(n4572), .ZN(n8909) );
  nd12d1 U4525 ( .A1(n17), .A2(n3009), .ZN(n8031) );
  nd04d1 U4526 ( .A1(n1342), .A2(n1299), .A3(n1247), .A4(n1563), .ZN(n17) );
  inv0d0 U4529 ( .I(n7620), .ZN(n4023) );
  nd02d1 U4530 ( .A1(n8857), .A2(n3798), .ZN(n5326) );
  inv0d0 U4531 ( .I(n5181), .ZN(n4318) );
  nd02d1 U4534 ( .A1(n3233), .A2(n3232), .ZN(n5562) );
  nr02d1 U4538 ( .A1(n6331), .A2(n5501), .ZN(n11766) );
  nd02d1 U4539 ( .A1(n11219), .A2(n11220), .ZN(n9438) );
  nd02d1 U4541 ( .A1(n11935), .A2(n4917), .ZN(n11939) );
  inv0d0 U4542 ( .I(n5712), .ZN(n5142) );
  nd02d1 U4543 ( .A1(n7392), .A2(n7393), .ZN(n7112) );
  nd02d1 U4544 ( .A1(N12450), .A2(n10837), .ZN(n9309) );
  nd03d1 U4547 ( .A1(n7444), .A2(n5458), .A3(n7562), .ZN(n8103) );
  inv0d0 U4550 ( .I(n7359), .ZN(n2998) );
  nd02d1 U4552 ( .A1(N9148), .A2(n8268), .ZN(n9777) );
  nd02d1 U4555 ( .A1(n7739), .A2(n3517), .ZN(n7748) );
  nd02d1 U4556 ( .A1(n5828), .A2(n5821), .ZN(n5020) );
  nd02d1 U4557 ( .A1(n5721), .A2(n7388), .ZN(n4981) );
  nd02d1 U4559 ( .A1(n3211), .A2(n3235), .ZN(n6416) );
  nd02d1 U4560 ( .A1(n9144), .A2(n3952), .ZN(n6632) );
  nd02d1 U4562 ( .A1(n5690), .A2(n4123), .ZN(n5908) );
  nd02d1 U4563 ( .A1(n3909), .A2(n3968), .ZN(n5117) );
  inv0d0 U4564 ( .I(n10126), .ZN(n3243) );
  nd02d1 U4566 ( .A1(N9036), .A2(n11416), .ZN(n11287) );
  nd03d1 U4567 ( .A1(n5364), .A2(n3224), .A3(N14050), .ZN(n6424) );
  nd02d1 U4569 ( .A1(N13970), .A2(n3235), .ZN(n8651) );
  nd03d1 U4571 ( .A1(n5096), .A2(n3944), .A3(N10446), .ZN(n7667) );
  nd02d1 U4574 ( .A1(N12386), .A2(n11681), .ZN(n5412) );
  nd02d1 U4575 ( .A1(n4008), .A2(n4013), .ZN(n5007) );
  nd02d1 U4577 ( .A1(n11839), .A2(n3084), .ZN(n4756) );
  inv0d0 U4578 ( .I(n4938), .ZN(n4998) );
  nd02d1 U4579 ( .A1(n3104), .A2(n3106), .ZN(n6499) );
  nd03d1 U4580 ( .A1(n6657), .A2(n5293), .A3(n11435), .ZN(n11439) );
  nr02d1 U4582 ( .A1(n6379), .A2(n3185), .ZN(n8634) );
  nr02d1 U4583 ( .A1(n6035), .A2(n5216), .ZN(n6036) );
  nd02d1 U4584 ( .A1(N11666), .A2(n12047), .ZN(n4446) );
  nd03d1 U4585 ( .A1(n4421), .A2(n5152), .A3(n3257), .ZN(n7178) );
  nd02d1 U4587 ( .A1(n4949), .A2(n8453), .ZN(n7015) );
  nd02d1 U4588 ( .A1(n5285), .A2(n4693), .ZN(n5294) );
  nr02d1 U4589 ( .A1(n6254), .A2(n6252), .ZN(n9355) );
  nd03d1 U4591 ( .A1(n3532), .A2(n3533), .A3(n3567), .ZN(n4449) );
  nd02d1 U4592 ( .A1(n5463), .A2(n5464), .ZN(n9369) );
  nr02d1 U4593 ( .A1(n5624), .A2(n5698), .ZN(n5638) );
  nr02d1 U4594 ( .A1(n6391), .A2(n7227), .ZN(n8637) );
  nd03d1 U4597 ( .A1(n6602), .A2(n4988), .A3(n7820), .ZN(n7827) );
  nr02d1 U4598 ( .A1(n5462), .A2(n3388), .ZN(n6263) );
  nd12d1 U4599 ( .A1(n18), .A2(n8147), .ZN(n8151) );
  nr04d1 U4600 ( .A1(n1182), .A2(n1138), .A3(n1239), .A4(n2669), .ZN(n18) );
  nr02d1 U4602 ( .A1(n9346), .A2(n9342), .ZN(n7823) );
  nd02d1 U4604 ( .A1(n2983), .A2(n2984), .ZN(n9538) );
  nd03d1 U4606 ( .A1(n4557), .A2(n4426), .A3(n4985), .ZN(n4562) );
  nr02d1 U4608 ( .A1(n9428), .A2(n6379), .ZN(n4664) );
  nr13d1 U4609 ( .A1(N10551), .A2(n8380), .A3(n6930), .ZN(n8383) );
  nr02d1 U4612 ( .A1(n2986), .A2(n10257), .ZN(n4830) );
  nd02d1 U4617 ( .A1(n4167), .A2(N9106), .ZN(n8110) );
  nd02d1 U4618 ( .A1(N15474), .A2(n2908), .ZN(n10327) );
  nd02d1 U4622 ( .A1(n7373), .A2(n4303), .ZN(n7249) );
  nd02d1 U4624 ( .A1(n10106), .A2(n7189), .ZN(n8066) );
  nr02d1 U4625 ( .A1(n4896), .A2(n4916), .ZN(n4903) );
  nd03d1 U4626 ( .A1(n5731), .A2(n5833), .A3(n7791), .ZN(n7798) );
  nr02d1 U4627 ( .A1(n4671), .A2(n3195), .ZN(n11985) );
  nd03d1 U4629 ( .A1(n4723), .A2(n4950), .A3(n5140), .ZN(n4740) );
  nd02d1 U4630 ( .A1(n5114), .A2(n5780), .ZN(n5127) );
  nd02d1 U4631 ( .A1(N11922), .A2(n3557), .ZN(n6143) );
  nd02d1 U4632 ( .A1(n8593), .A2(n8070), .ZN(n8597) );
  nd02d1 U4634 ( .A1(n7466), .A2(n4789), .ZN(n8144) );
  nd12d1 U4636 ( .A1(n19), .A2(n10257), .ZN(n10362) );
  nd04d1 U4639 ( .A1(n1342), .A2(n1300), .A3(n1246), .A4(n1520), .ZN(n19) );
  nd03d1 U4640 ( .A1(n3458), .A2(n3459), .A3(n11679), .ZN(n4508) );
  nd03d1 U4641 ( .A1(n4279), .A2(n9697), .A3(n5796), .ZN(n7496) );
  nd02d1 U4644 ( .A1(n4594), .A2(n4977), .ZN(n4605) );
  inv0d0 U4646 ( .I(n4896), .ZN(n2840) );
  oai211d1 U4649 ( .C1(n1230), .C2(n1279), .A(n1800), .B(n1337), .ZN(n20) );
  nr02d1 U4652 ( .A1(n2969), .A2(n4848), .ZN(n5662) );
  nd02d1 U4655 ( .A1(n6003), .A2(n3952), .ZN(n5177) );
  nd03d1 U4661 ( .A1(n4439), .A2(n3461), .A3(N12322), .ZN(n8526) );
  aoim22d1 U4666 ( .A1(n7274), .A2(n7275), .B1(n7276), .B2(n3055), .Z(n7273)
         );
  inv0d0 U4673 ( .I(n4737), .ZN(n3063) );
  nd02d1 U4676 ( .A1(N11890), .A2(n3559), .ZN(n5359) );
  nr02d1 U4685 ( .A1(n6188), .A2(n3362), .ZN(n7811) );
  nd02d1 U4687 ( .A1(n4595), .A2(n4628), .ZN(n7462) );
  nd02d1 U4695 ( .A1(N13314), .A2(n3283), .ZN(n11231) );
  nd02d1 U4696 ( .A1(N13186), .A2(n7160), .ZN(n7163) );
  nd02d1 U4701 ( .A1(n6134), .A2(n12047), .ZN(n12042) );
  nr02d1 U4710 ( .A1(n6643), .A2(n6644), .ZN(n6642) );
  inv0d0 U4730 ( .I(n5651), .ZN(n2965) );
  nd02d1 U4734 ( .A1(n3005), .A2(n3006), .ZN(n8043) );
  nd02d1 U4737 ( .A1(n5075), .A2(n7610), .ZN(n7617) );
  inv0d0 U4749 ( .I(n4826), .ZN(n2986) );
  inv0d0 U4754 ( .I(n7697), .ZN(n3848) );
  nd03d1 U4760 ( .A1(n5720), .A2(n3266), .A3(n3357), .ZN(n6286) );
  nd02d1 U4766 ( .A1(n7391), .A2(n3355), .ZN(n7119) );
  nd02d1 U4771 ( .A1(n6430), .A2(n9453), .ZN(n11010) );
  inv0d0 U4787 ( .I(n7557), .ZN(n4161) );
  nd03d1 U4789 ( .A1(n5380), .A2(n4972), .A3(n3265), .ZN(n11774) );
  nd03d1 U4794 ( .A1(n11430), .A2(n6139), .A3(N9204), .ZN(n5881) );
  nd03d1 U4796 ( .A1(n6663), .A2(n5693), .A3(n4747), .ZN(n5841) );
  nd02d1 U4799 ( .A1(n3065), .A2(n10384), .ZN(n5589) );
  nd02d1 U4801 ( .A1(n5837), .A2(n3793), .ZN(n11619) );
  inv0d0 U4813 ( .I(n5467), .ZN(n2807) );
  nd03d1 U4816 ( .A1(n4169), .A2(n5458), .A3(N9134), .ZN(n11283) );
  inv0d0 U4822 ( .I(n7078), .ZN(n3433) );
  nd02d1 U4828 ( .A1(n5237), .A2(n4714), .ZN(n4722) );
  nd02d1 U4829 ( .A1(n3038), .A2(n3128), .ZN(n10161) );
  nd02d1 U4831 ( .A1(n3076), .A2(n3077), .ZN(n11039) );
  inv0d0 U4834 ( .I(n5474), .ZN(n3273) );
  inv0d0 U4838 ( .I(n6030), .ZN(n3880) );
  nd03d1 U4842 ( .A1(n3838), .A2(n7685), .A3(N10746), .ZN(n9629) );
  nd02d1 U4844 ( .A1(n5406), .A2(n5833), .ZN(n4992) );
  nd03d1 U4845 ( .A1(n5271), .A2(n6117), .A3(n5261), .ZN(n5273) );
  nd02d1 U4846 ( .A1(n4991), .A2(n4529), .ZN(n4534) );
  nd02d1 U4851 ( .A1(n4055), .A2(n4742), .ZN(n11484) );
  nr02d1 U4857 ( .A1(n6379), .A2(n8626), .ZN(n7877) );
  nr23d1 U4858 ( .A1(n8005), .A2(n8006), .A3(n7340), .ZN(n8004) );
  nd02d1 U4860 ( .A1(n2993), .A2(n2994), .ZN(n7358) );
  nd02d1 U4865 ( .A1(n3546), .A2(n9255), .ZN(n5366) );
  nd02d1 U4866 ( .A1(n9563), .A2(n2876), .ZN(n9565) );
  nd02d1 U4868 ( .A1(n3889), .A2(n7421), .ZN(n7694) );
  nd02d1 U4875 ( .A1(N9711), .A2(n4055), .ZN(n11277) );
  nr02d1 U4876 ( .A1(n10812), .A2(n5382), .ZN(n9277) );
  nd03d1 U4883 ( .A1(n4985), .A2(n4426), .A3(n11711), .ZN(n11715) );
  nd03d1 U4886 ( .A1(n5237), .A2(n5729), .A3(n5572), .ZN(n5576) );
  nd03d1 U4887 ( .A1(n12059), .A2(n3821), .A3(N10596), .ZN(n11556) );
  nd02d1 U4894 ( .A1(n6787), .A2(n4071), .ZN(n5032) );
  inv0d0 U4898 ( .I(n6028), .ZN(n3879) );
  nd02d1 U4909 ( .A1(n3928), .A2(n8356), .ZN(n4422) );
  inv0d0 U4910 ( .I(n5375), .ZN(n3479) );
  nd03d1 U4917 ( .A1(n3913), .A2(n3968), .A3(n5120), .ZN(n7653) );
  nd03d1 U4923 ( .A1(n4303), .A2(n4960), .A3(n11808), .ZN(n11815) );
  nd03d1 U4928 ( .A1(n4985), .A2(n5724), .A3(n3359), .ZN(n6239) );
  nd02d1 U4931 ( .A1(n5719), .A2(n10106), .ZN(n8606) );
  nr02d1 U4932 ( .A1(n3152), .A2(n5142), .ZN(n8633) );
  nd03d1 U4938 ( .A1(n3802), .A2(n5939), .A3(N11346), .ZN(n10732) );
  nd02d1 U4963 ( .A1(n5331), .A2(n3787), .ZN(n6109) );
  inv0d0 U4965 ( .I(n6593), .ZN(n3297) );
  nd02d1 U4968 ( .A1(N11541), .A2(n11622), .ZN(n6122) );
  nd02d1 U4969 ( .A1(n11395), .A2(n5697), .ZN(n11402) );
  nr02d1 U4972 ( .A1(n7628), .A2(n8094), .ZN(n7636) );
  nd03d1 U4975 ( .A1(n8862), .A2(n3870), .A3(N10971), .ZN(n6961) );
  inv0d0 U4982 ( .I(n6169), .ZN(n3472) );
  nd03d1 U4984 ( .A1(n3503), .A2(n5414), .A3(n4944), .ZN(n7774) );
  nd02d1 U4989 ( .A1(n8026), .A2(n2904), .ZN(n8016) );
  inv0d0 U4990 ( .I(n4729), .ZN(n3127) );
  nd02d1 U4991 ( .A1(n4895), .A2(n3013), .ZN(n7972) );
  inv0d0 U4992 ( .I(n6258), .ZN(n3398) );
  nd02d1 U4993 ( .A1(n8988), .A2(n4205), .ZN(n11385) );
  inv0d0 U4995 ( .I(n8283), .ZN(n4127) );
  nd03d1 U4996 ( .A1(n4481), .A2(n5783), .A3(n5441), .ZN(n5107) );
  nd02d1 U4997 ( .A1(n7135), .A2(n11720), .ZN(n4565) );
  nd02d1 U4999 ( .A1(n4229), .A2(n7455), .ZN(n11366) );
  nd02d1 U5001 ( .A1(n3186), .A2(n3187), .ZN(n9428) );
  nr02d1 U5004 ( .A1(n10493), .A2(n12072), .ZN(n11357) );
  nd03d1 U5005 ( .A1(n4152), .A2(n4154), .A3(n5828), .ZN(n5823) );
  inv0d0 U5006 ( .I(n10245), .ZN(n2917) );
  nd02d1 U5007 ( .A1(n5367), .A2(n10788), .ZN(n10003) );
  nd03d1 U5013 ( .A1(n4239), .A2(n8119), .A3(N8406), .ZN(n11348) );
  nd03d1 U5014 ( .A1(n3921), .A2(n3964), .A3(N10221), .ZN(n5137) );
  inv0d0 U5020 ( .I(n10863), .ZN(n3416) );
  nd12d1 U5021 ( .A1(n21), .A2(n4819), .ZN(n8146) );
  nr04d1 U5023 ( .A1(n1341), .A2(n1295), .A3(n1239), .A4(n2673), .ZN(n21) );
  nd02d1 U5025 ( .A1(n3222), .A2(n3220), .ZN(n8661) );
  nd02d1 U5026 ( .A1(N10176), .A2(n3966), .ZN(n9860) );
  nd02d1 U5028 ( .A1(n5720), .A2(n9370), .ZN(n9377) );
  inv0d0 U5029 ( .I(n6154), .ZN(n3551) );
  nd02d1 U5030 ( .A1(n4814), .A2(n7336), .ZN(n4815) );
  nd02d1 U5031 ( .A1(n2910), .A2(n2911), .ZN(n11140) );
  nd02d1 U5032 ( .A1(n4576), .A2(n4561), .ZN(n8919) );
  nd02d1 U5033 ( .A1(n3548), .A2(n10788), .ZN(n9617) );
  nd02d1 U5034 ( .A1(n8866), .A2(n3963), .ZN(n5153) );
  nd02d1 U5036 ( .A1(n3872), .A2(n3870), .ZN(n7417) );
  nd02d1 U5037 ( .A1(n11687), .A2(n4991), .ZN(n11693) );
  nd02d1 U5043 ( .A1(n3017), .A2(n3105), .ZN(n9491) );
  nd02d1 U5045 ( .A1(n3017), .A2(n6500), .ZN(n4774) );
  nd02d1 U5046 ( .A1(N10506), .A2(n10657), .ZN(n10661) );
  nd02d1 U5049 ( .A1(n5435), .A2(n10657), .ZN(n5180) );
  nd02d1 U5053 ( .A1(N10086), .A2(n4044), .ZN(n5976) );
  nd02d1 U5054 ( .A1(N14354), .A2(n3077), .ZN(n8707) );
  inv0d0 U5060 ( .I(n1610), .ZN(n1613) );
  nd02d1 U5062 ( .A1(n7660), .A2(n5093), .ZN(n7661) );
  nd02d1 U5063 ( .A1(n4290), .A2(n7453), .ZN(n8113) );
  nd02d1 U5064 ( .A1(n5188), .A2(n5767), .ZN(n5196) );
  inv0d0 U5065 ( .I(n6301), .ZN(n3321) );
  nd02d1 U5069 ( .A1(n3496), .A2(n4996), .ZN(n11667) );
  nd02d1 U5070 ( .A1(n3502), .A2(n4996), .ZN(n4499) );
  nd02d1 U5072 ( .A1(n7122), .A2(n5634), .ZN(n7126) );
  nd03d1 U5074 ( .A1(n4019), .A2(n12063), .A3(N9801), .ZN(n8322) );
  nd12d1 U5076 ( .A1(n22), .A2(n2886), .ZN(n10322) );
  nd04d1 U5077 ( .A1(n1304), .A2(n1244), .A3(n1340), .A4(n1453), .ZN(n22) );
  nd02d1 U5078 ( .A1(N10251), .A2(n3963), .ZN(n6893) );
  nd02d1 U5079 ( .A1(n4113), .A2(n6657), .ZN(n5899) );
  inv0d0 U5080 ( .I(n7409), .ZN(n4683) );
  nd02d1 U5081 ( .A1(n3238), .A2(n3239), .ZN(n6407) );
  inv0d0 U5082 ( .I(n5464), .ZN(n3391) );
  nd03d1 U5083 ( .A1(n5071), .A2(n3873), .A3(N10926), .ZN(n5244) );
  nd02d1 U5084 ( .A1(n3288), .A2(n3286), .ZN(n6320) );
  inv0d0 U5087 ( .I(n7392), .ZN(n3487) );
  inv0d0 U5091 ( .I(n8836), .ZN(n3240) );
  nd02d1 U5092 ( .A1(n11625), .A2(n5345), .ZN(n11627) );
  nd02d1 U5095 ( .A1(N10641), .A2(n6013), .ZN(n6022) );
  nd02d1 U5096 ( .A1(n5165), .A2(n3467), .ZN(n5395) );
  nd02d1 U5097 ( .A1(n6018), .A2(n7064), .ZN(n8507) );
  nd02d1 U5099 ( .A1(N13170), .A2(n11741), .ZN(n11738) );
  nd02d1 U5105 ( .A1(n3965), .A2(n4725), .ZN(n7652) );
  nd03d1 U5110 ( .A1(n4977), .A2(n5152), .A3(n6302), .ZN(n6307) );
  inv0d0 U5111 ( .I(n10500), .ZN(n4269) );
  nd02d1 U5112 ( .A1(n2925), .A2(n4790), .ZN(n5628) );
  nd02d1 U5113 ( .A1(n3239), .A2(n3235), .ZN(n8649) );
  nd03d1 U5116 ( .A1(n6652), .A2(n5579), .A3(n11454), .ZN(n11462) );
  nd02d1 U5117 ( .A1(n4153), .A2(n4152), .ZN(n5039) );
  nd02d1 U5118 ( .A1(n8486), .A2(n9998), .ZN(n7041) );
  nd02d1 U5120 ( .A1(n4810), .A2(n4822), .ZN(n6522) );
  nd12d1 U5121 ( .A1(n2298), .A2(n7648), .ZN(n7650) );
  nd03d1 U5122 ( .A1(n5693), .A2(n6665), .A3(n4214), .ZN(n6754) );
  nd02d1 U5128 ( .A1(N11938), .A2(n3546), .ZN(n5363) );
  nd02d1 U5129 ( .A1(n4063), .A2(n5888), .ZN(n5884) );
  nd02d1 U5132 ( .A1(N10326), .A2(n6902), .ZN(n10640) );
  nd02d1 U5133 ( .A1(n7003), .A2(n11615), .ZN(n9221) );
  nd02d1 U5135 ( .A1(n8069), .A2(n3285), .ZN(n4615) );
  nd02d1 U5136 ( .A1(n4036), .A2(n4034), .ZN(n7437) );
  inv0d0 U5137 ( .I(n10384), .ZN(n3122) );
  nd02d1 U5138 ( .A1(n8785), .A2(n2983), .ZN(n10271) );
  nd12d1 U5140 ( .A1(n23), .A2(n2993), .ZN(n11873) );
  nd04d1 U5141 ( .A1(n1342), .A2(n1300), .A3(n1534), .A4(n1242), .ZN(n23) );
  nd02d1 U5142 ( .A1(n4784), .A2(n5224), .ZN(n4801) );
  nd02d1 U5144 ( .A1(n3740), .A2(n3748), .ZN(n9940) );
  nd02d1 U5145 ( .A1(N8342), .A2(n11338), .ZN(n9696) );
  nd02d1 U5147 ( .A1(n3865), .A2(n3858), .ZN(n8423) );
  nd03d1 U5148 ( .A1(n6623), .A2(n5271), .A3(n3883), .ZN(n11588) );
  inv0d0 U5149 ( .I(n10013), .ZN(n3473) );
  nd02d1 U5150 ( .A1(N8186), .A2(n4572), .ZN(n9670) );
  nd02d1 U5151 ( .A1(N9786), .A2(n4020), .ZN(n8321) );
  nd02d1 U5152 ( .A1(N9414), .A2(n12064), .ZN(n8297) );
  nd02d1 U5154 ( .A1(n3969), .A2(n7647), .ZN(n5115) );
  nd02d1 U5157 ( .A1(n5783), .A2(n5101), .ZN(n8094) );
  nd03d1 U5158 ( .A1(n4013), .A2(n8317), .A3(n6648), .ZN(n5965) );
  nd02d1 U5159 ( .A1(n3801), .A2(n3774), .ZN(n6094) );
  nd02d1 U5160 ( .A1(n4792), .A2(n3007), .ZN(n4795) );
  nd02d1 U5162 ( .A1(n5344), .A2(n6561), .ZN(n5699) );
  nd02d1 U5165 ( .A1(n3799), .A2(n10407), .ZN(n10735) );
  nr02d1 U5166 ( .A1(n6616), .A2(n4456), .ZN(n9250) );
  nd02d1 U5168 ( .A1(N9232), .A2(n5888), .ZN(n7569) );
  nd02d1 U5169 ( .A1(n3876), .A2(n5550), .ZN(n5239) );
  nd02d1 U5170 ( .A1(n7922), .A2(n3044), .ZN(n8672) );
  nr02d1 U5173 ( .A1(n7755), .A2(n8076), .ZN(n7758) );
  nd02d1 U5174 ( .A1(N9386), .A2(n4080), .ZN(n5915) );
  nd02d1 U5175 ( .A1(N9022), .A2(n9018), .ZN(n10544) );
  nd02d1 U5176 ( .A1(n11336), .A2(n8126), .ZN(n10472) );
  nd02d1 U5178 ( .A1(n8867), .A2(n3920), .ZN(n5132) );
  nd02d1 U5181 ( .A1(n11605), .A2(n5182), .ZN(n5305) );
  nd02d1 U5183 ( .A1(n7040), .A2(n3561), .ZN(n6615) );
  nd02d1 U5185 ( .A1(n4111), .A2(n5909), .ZN(n9791) );
  nd02d1 U5186 ( .A1(n5124), .A2(n11932), .ZN(n11142) );
  nd02d1 U5190 ( .A1(n3950), .A2(n9144), .ZN(n5773) );
  nd02d1 U5193 ( .A1(N11016), .A2(n11583), .ZN(n9929) );
  nd02d1 U5199 ( .A1(N9316), .A2(n8282), .ZN(n6791) );
  nd02d1 U5200 ( .A1(n10825), .A2(n3466), .ZN(n9294) );
  nr02d1 U5204 ( .A1(n9315), .A2(n6194), .ZN(n7804) );
  nd02d1 U5207 ( .A1(n5914), .A2(n4075), .ZN(n6803) );
  nd03d1 U5210 ( .A1(n3252), .A2(n4972), .A3(n5380), .ZN(n4632) );
  nd02d1 U5219 ( .A1(n2896), .A2(n11175), .ZN(n10339) );
  inv0d0 U5228 ( .I(n5717), .ZN(n4423) );
  inv0d0 U5230 ( .I(n8116), .ZN(n4264) );
  nd02d1 U5236 ( .A1(N12706), .A2(n12017), .ZN(n9336) );
  inv0d0 U5237 ( .I(n1870), .ZN(N12706) );
  inv0d0 U5247 ( .I(n1869), .ZN(n1871) );
  nd02d1 U5248 ( .A1(n3168), .A2(n3167), .ZN(n10120) );
  nd02d1 U5250 ( .A1(n8266), .A2(n5872), .ZN(n5037) );
  nd02d1 U5253 ( .A1(n6973), .A2(n4692), .ZN(n6980) );
  inv0d0 U5261 ( .I(n7100), .ZN(n3453) );
  inv0d0 U5267 ( .I(n7088), .ZN(n3488) );
  nd03d1 U5270 ( .A1(n5380), .A2(n4972), .A3(n3267), .ZN(n7871) );
  inv0d0 U5279 ( .I(n7333), .ZN(n2974) );
  nd02d1 U5296 ( .A1(n5724), .A2(n6602), .ZN(n12003) );
  inv0d0 U5297 ( .I(n11478), .ZN(n3994) );
  nd03d1 U5304 ( .A1(n11219), .A2(n3239), .A3(n3208), .ZN(n8059) );
  nd03d1 U5305 ( .A1(n5529), .A2(n3204), .A3(n3238), .ZN(n7241) );
  nd02d1 U5307 ( .A1(n2992), .A2(n11971), .ZN(n10369) );
  nd02d1 U5309 ( .A1(n4228), .A2(n7453), .ZN(n11384) );
  nd03d1 U5311 ( .A1(n5752), .A2(n4457), .A3(n6078), .ZN(n6091) );
  inv0d0 U5312 ( .I(n8153), .ZN(n4523) );
  nd03d1 U5313 ( .A1(n5751), .A2(n5752), .A3(n3665), .ZN(n11610) );
  inv0d0 U5316 ( .I(n5529), .ZN(n3197) );
  nd02d1 U5317 ( .A1(N12690), .A2(n12016), .ZN(n10869) );
  nd02d1 U5320 ( .A1(n4457), .A2(n3804), .ZN(n10728) );
  nd02d1 U5325 ( .A1(N10866), .A2(n3876), .ZN(n6951) );
  nd02d1 U5327 ( .A1(n5424), .A2(n3446), .ZN(n8547) );
  nd02d1 U5330 ( .A1(n7987), .A2(n4842), .ZN(n6536) );
  inv0d0 U5339 ( .I(n5222), .ZN(n3897) );
  nr02d1 U5344 ( .A1(n7236), .A2(n8642), .ZN(n10142) );
  inv0d0 U5351 ( .I(n7511), .ZN(n4255) );
  nd02d1 U5357 ( .A1(n5529), .A2(n7227), .ZN(n7893) );
  inv0d0 U5360 ( .I(n8920), .ZN(n4530) );
  inv0d0 U5361 ( .I(n9310), .ZN(n3454) );
  nd02d1 U5362 ( .A1(n8483), .A2(n4444), .ZN(n8481) );
  inv0d0 U5365 ( .I(n6635), .ZN(n3974) );
  nd02d1 U5381 ( .A1(n5120), .A2(n3967), .ZN(n5781) );
  inv0d0 U5383 ( .I(n6824), .ZN(n4133) );
  nr13d1 U5390 ( .A1(n4977), .A2(n4978), .A3(n5472), .ZN(n5481) );
  inv0d0 U5392 ( .I(n7235), .ZN(n3193) );
  inv0d0 U5395 ( .I(n8827), .ZN(n2895) );
  nd02d1 U5403 ( .A1(n11629), .A2(n4442), .ZN(n11633) );
  nd03d1 U5410 ( .A1(n2828), .A2(n7335), .A3(n6549), .ZN(n4931) );
  nd02d1 U5412 ( .A1(n7633), .A2(n10617), .ZN(n6644) );
  inv0d0 U5413 ( .I(n5331), .ZN(n3781) );
  inv0d0 U5420 ( .I(n8076), .ZN(n4444) );
  nd02d1 U5423 ( .A1(N10191), .A2(n3965), .ZN(n5131) );
  inv0d0 U5435 ( .I(n2278), .ZN(n2281) );
  inv0d0 U5437 ( .I(n8341), .ZN(n3907) );
  nd03d1 U5439 ( .A1(n3023), .A2(n5904), .A3(n4411), .ZN(n4750) );
  nd02d1 U5442 ( .A1(N12338), .A2(n3439), .ZN(n11672) );
  nd02d1 U5445 ( .A1(N13874), .A2(n3200), .ZN(n7890) );
  nd02d1 U5457 ( .A1(N10401), .A2(n6910), .ZN(n6913) );
  nd02d1 U5461 ( .A1(n8383), .A2(n12059), .ZN(n12060) );
  nd02d1 U5465 ( .A1(n4183), .A2(n9008), .ZN(n9004) );
  nd02d1 U5468 ( .A1(n4684), .A2(n4960), .ZN(n4688) );
  nd02d1 U5470 ( .A1(N10566), .A2(n12059), .ZN(n10663) );
  nd02d1 U5471 ( .A1(n3788), .A2(n11622), .ZN(n11626) );
  nd03d1 U5480 ( .A1(n4962), .A2(n5441), .A3(n7636), .ZN(n7642) );
  nd02d1 U5481 ( .A1(n6227), .A2(n4988), .ZN(n6222) );
  nd03d1 U5486 ( .A1(n4199), .A2(n5779), .A3(N8784), .ZN(n9737) );
  nd02d1 U5490 ( .A1(N13122), .A2(n12002), .ZN(n10910) );
  nd02d1 U5492 ( .A1(N8718), .A2(n8988), .ZN(n8986) );
  nd02d1 U5493 ( .A1(n3439), .A2(n3460), .ZN(n7401) );
  nd02d1 U5496 ( .A1(n7932), .A2(n4730), .ZN(n7936) );
  inv0d0 U5512 ( .I(n6252), .ZN(n3399) );
  nd02d1 U5513 ( .A1(n11736), .A2(n4656), .ZN(n11743) );
  nd02d1 U5519 ( .A1(n4405), .A2(n5129), .ZN(n6551) );
  nd02d1 U5523 ( .A1(N10386), .A2(n3938), .ZN(n11540) );
  nd02d1 U5525 ( .A1(n5469), .A2(n5720), .ZN(n5472) );
  nr02d1 U5527 ( .A1(n8627), .A2(n10126), .ZN(n4659) );
  nd02d1 U5535 ( .A1(n4656), .A2(n5252), .ZN(n4978) );
  nr02d1 U5540 ( .A1(n6694), .A2(n4277), .ZN(n11344) );
  nd02d1 U5547 ( .A1(n4683), .A2(n6134), .ZN(n5004) );
  nd02d1 U5549 ( .A1(N13330), .A2(n11753), .ZN(n11229) );
  nd03d1 U5551 ( .A1(n4510), .A2(n6663), .A3(n4213), .ZN(n6755) );
  nd02d1 U5552 ( .A1(n7903), .A2(n4960), .ZN(n7905) );
  inv0d0 U5553 ( .I(n9807), .ZN(n4059) );
  inv0d0 U5554 ( .I(n7373), .ZN(n3144) );
  nd02d1 U5556 ( .A1(n6514), .A2(n4940), .ZN(n6518) );
  inv0d0 U5558 ( .I(n4529), .ZN(n3501) );
  inv0d0 U5559 ( .I(n12026), .ZN(n3556) );
  nd02d1 U5561 ( .A1(n6883), .A2(n3921), .ZN(n6878) );
  inv0d0 U5564 ( .I(n8957), .ZN(n4271) );
  nd02d1 U5567 ( .A1(N8510), .A2(n4250), .ZN(n8954) );
  nd02d1 U5568 ( .A1(n4247), .A2(n8197), .ZN(n10491) );
  nd03d1 U5570 ( .A1(n5690), .A2(n6656), .A3(n4138), .ZN(n11448) );
  nd02d1 U5572 ( .A1(n5592), .A2(n4411), .ZN(n5596) );
  nd03d1 U5573 ( .A1(n5642), .A2(n6018), .A3(n7061), .ZN(n7070) );
  inv0d0 U5576 ( .I(n6003), .ZN(n3946) );
  nd03d1 U5577 ( .A1(n3972), .A2(n5683), .A3(n6045), .ZN(n5148) );
  nd03d1 U5578 ( .A1(n5427), .A2(n5837), .A3(n5327), .ZN(n5335) );
  nd02d1 U5579 ( .A1(n3148), .A2(n5711), .ZN(n11802) );
  nd03d1 U5580 ( .A1(n5101), .A2(n5570), .A3(n11498), .ZN(n11504) );
  nd02d1 U5581 ( .A1(N15250), .A2(n2864), .ZN(n9590) );
  nd03d1 U5582 ( .A1(n4913), .A2(n3146), .A3(n5508), .ZN(n5511) );
  inv0d0 U5584 ( .I(n9500), .ZN(n3011) );
  inv0d0 U5586 ( .I(n11220), .ZN(n3206) );
  inv0d0 U5587 ( .I(n7675), .ZN(n3834) );
  nd02d1 U5589 ( .A1(n3309), .A2(n10106), .ZN(n9402) );
  nd02d1 U5591 ( .A1(n3826), .A2(n6013), .ZN(n6941) );
  nd02d1 U5592 ( .A1(N12290), .A2(n3461), .ZN(n10828) );
  nd02d1 U5594 ( .A1(N9176), .A2(n11430), .ZN(n9776) );
  nr02d1 U5595 ( .A1(n7831), .A2(n12003), .ZN(n4987) );
  nd03d1 U5596 ( .A1(n5852), .A2(n5582), .A3(n4207), .ZN(n7559) );
  inv0d0 U5597 ( .I(n5042), .ZN(n4155) );
  nd02d1 U5598 ( .A1(N12114), .A2(n3475), .ZN(n10812) );
  inv0d0 U5599 ( .I(n1964), .ZN(N12114) );
  inv0d0 U5601 ( .I(n7548), .ZN(n4177) );
  nd02d1 U5603 ( .A1(n3939), .A2(n3943), .ZN(n5999) );
  nd02d1 U5604 ( .A1(n4272), .A2(n4273), .ZN(n10493) );
  nd02d1 U5605 ( .A1(n4181), .A2(n6663), .ZN(n7539) );
  nd03d1 U5606 ( .A1(n3218), .A2(n4901), .A3(n7252), .ZN(n7256) );
  nd02d1 U5607 ( .A1(n5734), .A2(n7112), .ZN(n7114) );
  nd03d1 U5608 ( .A1(n3770), .A2(n3800), .A3(n3773), .ZN(n9954) );
  inv0d0 U5613 ( .I(n5865), .ZN(n4324) );
  inv0d0 U5616 ( .I(n11338), .ZN(n4277) );
  nd02d1 U5617 ( .A1(n5987), .A2(n3159), .ZN(n4657) );
  inv0d0 U5618 ( .I(n7463), .ZN(n4771) );
  inv0d0 U5619 ( .I(n7838), .ZN(n3384) );
  nd02d1 U5620 ( .A1(n3326), .A2(n7160), .ZN(n7161) );
  nd03d1 U5624 ( .A1(n7751), .A2(n3526), .A3(n3569), .ZN(n6130) );
  inv0d0 U5627 ( .I(n8642), .ZN(n3192) );
  inv0d0 U5630 ( .I(n6114), .ZN(n3681) );
  inv0d0 U5632 ( .I(n11721), .ZN(n3395) );
  nd02d1 U5634 ( .A1(n8580), .A2(n3266), .ZN(n8584) );
  nd02d1 U5636 ( .A1(n5152), .A2(n6311), .ZN(n7175) );
  nd02d1 U5638 ( .A1(n4108), .A2(n4106), .ZN(n5923) );
  nd03d1 U5640 ( .A1(n3158), .A2(n5364), .A3(n4901), .ZN(n4697) );
  nd02d1 U5643 ( .A1(n8413), .A2(n3875), .ZN(n9919) );
  nd02d1 U5644 ( .A1(N8162), .A2(n4590), .ZN(n11323) );
  nd02d1 U5645 ( .A1(n3981), .A2(n6888), .ZN(n9128) );
  nd02d1 U5646 ( .A1(n5274), .A2(n4693), .ZN(n8081) );
  nd03d1 U5647 ( .A1(n4066), .A2(n11439), .A3(n5895), .ZN(n11438) );
  inv0d0 U5649 ( .I(n5874), .ZN(n4117) );
  inv0d0 U5653 ( .I(n5491), .ZN(n3291) );
  inv0d0 U5654 ( .I(n7223), .ZN(n3244) );
  nd02d1 U5656 ( .A1(n4767), .A2(n8131), .ZN(n10441) );
  inv0d0 U5659 ( .I(n9239), .ZN(n3569) );
  nd02d1 U5661 ( .A1(N9246), .A2(n4115), .ZN(n10555) );
  inv0d0 U5662 ( .I(n11677), .ZN(n5535) );
  inv0d0 U5663 ( .I(n9816), .ZN(n3985) );
  nd02d1 U5664 ( .A1(n4201), .A2(n5778), .ZN(n8995) );
  nd02d1 U5665 ( .A1(n4693), .A2(n9199), .ZN(n9939) );
  nd12d1 U5666 ( .A1(n2654), .A2(n4392), .ZN(n8922) );
  nd02d1 U5670 ( .A1(N9981), .A2(n4048), .ZN(n9839) );
  nd02d1 U5672 ( .A1(N8367), .A2(n11342), .ZN(n6690) );
  inv0d0 U5674 ( .I(n2625), .ZN(N8367) );
  nd02d1 U5675 ( .A1(n3035), .A2(n3128), .ZN(n7915) );
  nd02d1 U5678 ( .A1(n7864), .A2(n5044), .ZN(n7867) );
  inv0d0 U5680 ( .I(n6194), .ZN(n3444) );
  nd02d1 U5681 ( .A1(n4184), .A2(n6665), .ZN(n8241) );
  nd02d1 U5682 ( .A1(n11757), .A2(n5044), .ZN(n11762) );
  nd02d1 U5683 ( .A1(n4869), .A2(n10288), .ZN(n9594) );
  nd02d1 U5684 ( .A1(n4078), .A2(n4108), .ZN(n9795) );
  nd02d1 U5685 ( .A1(n4175), .A2(n11416), .ZN(n9761) );
  nd02d1 U5688 ( .A1(n4180), .A2(n4510), .ZN(n11409) );
  nd02d1 U5694 ( .A1(n11896), .A2(n4927), .ZN(n11899) );
  nd02d1 U5695 ( .A1(n5674), .A2(n4927), .ZN(n5677) );
  nd02d1 U5696 ( .A1(N14658), .A2(n3010), .ZN(n11853) );
  inv0d0 U5697 ( .I(n7258), .ZN(n3229) );
  nd02d1 U5698 ( .A1(n3084), .A2(n3116), .ZN(n9602) );
  nd02d1 U5702 ( .A1(n7450), .A2(n4510), .ZN(n5844) );
  nd02d1 U5703 ( .A1(n11951), .A2(n4910), .ZN(n11952) );
  nd03d1 U5704 ( .A1(n6623), .A2(n4954), .A3(n3888), .ZN(n7709) );
  nd03d1 U5706 ( .A1(n4901), .A2(n5364), .A3(n3155), .ZN(n7912) );
  inv0d0 U5709 ( .I(n5706), .ZN(n3024) );
  nd02d1 U5710 ( .A1(n10935), .A2(n3288), .ZN(n10102) );
  nd02d1 U5712 ( .A1(n4369), .A2(n4357), .ZN(n6679) );
  nd02d1 U5715 ( .A1(n6044), .A2(n5759), .ZN(n6047) );
  inv0d0 U5717 ( .I(n10025), .ZN(n3483) );
  inv0d0 U5720 ( .I(n7226), .ZN(n3143) );
  nd02d1 U5723 ( .A1(n4927), .A2(n4853), .ZN(n4861) );
  nd02d1 U5726 ( .A1(n6656), .A2(n4124), .ZN(n5901) );
  inv0d0 U5727 ( .I(n5399), .ZN(n3481) );
  nd02d1 U5729 ( .A1(n3472), .A2(n6167), .ZN(n9285) );
  nd02d1 U5730 ( .A1(n7217), .A2(n3249), .ZN(n10963) );
  nd02d1 U5731 ( .A1(n3840), .A2(n3878), .ZN(n5215) );
  nd02d1 U5732 ( .A1(n11589), .A2(n5748), .ZN(n11592) );
  nd02d1 U5733 ( .A1(n5101), .A2(n4051), .ZN(n7631) );
  nd02d1 U5736 ( .A1(n4052), .A2(n5570), .ZN(n5087) );
  inv0d0 U5739 ( .I(n6899), .ZN(n3928) );
  inv0d0 U5740 ( .I(n6364), .ZN(n3249) );
  nd02d1 U5741 ( .A1(n5044), .A2(n4612), .ZN(n4625) );
  inv0d0 U5745 ( .I(n8369), .ZN(n3983) );
  inv0d0 U5747 ( .I(n4814), .ZN(n3002) );
  nd02d1 U5748 ( .A1(N10416), .A2(n3944), .ZN(n10648) );
  nd03d1 U5749 ( .A1(n4922), .A2(n5389), .A3(n7832), .ZN(n7842) );
  nd02d1 U5753 ( .A1(N11211), .A2(n3807), .ZN(n5297) );
  nd02d1 U5754 ( .A1(n3010), .A2(n2926), .ZN(n4783) );
  nd02d1 U5755 ( .A1(n4683), .A2(n6124), .ZN(n6129) );
  inv0d0 U5756 ( .I(n10892), .ZN(n3397) );
  nd02d1 U5759 ( .A1(n4312), .A2(n3559), .ZN(n6145) );
  inv0d0 U5760 ( .I(n9342), .ZN(n3404) );
  nd02d1 U5761 ( .A1(N13138), .A2(n12001), .ZN(n10912) );
  nd02d1 U5764 ( .A1(N15330), .A2(n11932), .ZN(n11189) );
  nd02d1 U5772 ( .A1(n5693), .A2(n4182), .ZN(n6757) );
  nd02d1 U5773 ( .A1(n3668), .A2(n6033), .ZN(n11601) );
  nd02d1 U5774 ( .A1(N10491), .A2(n3953), .ZN(n11549) );
  inv0d0 U5775 ( .I(n6985), .ZN(n3761) );
  inv0d0 U5776 ( .I(n10288), .ZN(n2852) );
  inv0d0 U5784 ( .I(n11703), .ZN(n3347) );
  nd02d1 U5789 ( .A1(n3882), .A2(n3826), .ZN(n9896) );
  nd02d1 U5793 ( .A1(N10656), .A2(n3835), .ZN(n6942) );
  inv0d0 U5808 ( .I(n8483), .ZN(n3515) );
  nd02d1 U5813 ( .A1(N8210), .A2(n11324), .ZN(n10463) );
  nd02d1 U5818 ( .A1(n2835), .A2(n4925), .ZN(n11914) );
  inv0d0 U5821 ( .I(n11770), .ZN(n3312) );
  nd02d1 U5826 ( .A1(n3856), .A2(n3854), .ZN(n7700) );
  nd02d1 U5827 ( .A1(n3421), .A2(n6198), .ZN(n8854) );
  inv0d0 U5830 ( .I(n8869), .ZN(n3982) );
  nd02d1 U5833 ( .A1(n6269), .A2(n4922), .ZN(n6274) );
  nd02d1 U5835 ( .A1(n3401), .A2(n6232), .ZN(n10077) );
  inv0d0 U5844 ( .I(n4478), .ZN(n3424) );
  nd02d1 U5845 ( .A1(n8839), .A2(n6593), .ZN(n8845) );
  nd02d1 U5850 ( .A1(n3973), .A2(n4711), .ZN(n5149) );
  nd02d1 U5856 ( .A1(n5331), .A2(n11619), .ZN(n7743) );
  inv0d0 U5857 ( .I(n4559), .ZN(n3378) );
  inv0d0 U5860 ( .I(n10057), .ZN(n3366) );
  inv0d0 U5863 ( .I(n7418), .ZN(n3868) );
  nd02d1 U5868 ( .A1(n5088), .A2(n4050), .ZN(n5975) );
  nd03d1 U5869 ( .A1(n4962), .A2(n8869), .A3(n8336), .ZN(n8346) );
  nd02d1 U5870 ( .A1(n2882), .A2(n2876), .ZN(n11928) );
  nd02d1 U5873 ( .A1(n3344), .A2(n6602), .ZN(n9349) );
  nd02d1 U5874 ( .A1(n7691), .A2(n5219), .ZN(n6043) );
  inv0d0 U5885 ( .I(n7760), .ZN(n3538) );
  inv0d0 U5886 ( .I(n11430), .ZN(n4061) );
  inv0d0 U5888 ( .I(n5745), .ZN(n3564) );
  nd03d1 U5892 ( .A1(n3956), .A2(n11556), .A3(n3817), .ZN(n9892) );
  nd02d1 U5903 ( .A1(n4956), .A2(n4701), .ZN(n4712) );
  nd02d1 U5904 ( .A1(n7145), .A2(n3266), .ZN(n7146) );
  inv0d0 U5906 ( .I(n8356), .ZN(n3926) );
  inv0d0 U5907 ( .I(n8389), .ZN(n3894) );
  inv0d0 U5910 ( .I(n7025), .ZN(n3517) );
  inv0d0 U5912 ( .I(n8549), .ZN(n3418) );
  inv0d0 U5913 ( .I(n5448), .ZN(n3335) );
  inv0d0 U5916 ( .I(n5501), .ZN(n3309) );
  nd02d1 U5917 ( .A1(n5751), .A2(n5304), .ZN(n5316) );
  inv0d0 U5922 ( .I(n5016), .ZN(n4163) );
  inv0d0 U5925 ( .I(n6835), .ZN(n4097) );
  inv0d0 U5926 ( .I(n9092), .ZN(n3990) );
  inv0d0 U5928 ( .I(n8246), .ZN(n4220) );
  inv0d0 U5929 ( .I(n11622), .ZN(n3522) );
  nd02d1 U5936 ( .A1(n11450), .A2(n7440), .ZN(n11457) );
  inv0d0 U5937 ( .I(n5637), .ZN(n2942) );
  inv0d0 U5940 ( .I(n6517), .ZN(n2954) );
  inv0d0 U5941 ( .I(n5403), .ZN(n3435) );
  nd02d1 U5944 ( .A1(n8668), .A2(n5706), .ZN(n8678) );
  inv0d0 U5951 ( .I(n10444), .ZN(n4881) );
  inv0d0 U5960 ( .I(n9895), .ZN(n3812) );
  inv0d0 U5961 ( .I(n7919), .ZN(n3038) );
  inv0d0 U5965 ( .I(n7002), .ZN(n3795) );
  inv0d0 U5972 ( .I(n11961), .ZN(n2855) );
  nd03d1 U5974 ( .A1(n4438), .A2(n5642), .A3(n7782), .ZN(n7784) );
  inv0d0 U5975 ( .I(n9037), .ZN(n4139) );
  inv0d1 U5980 ( .I(n1030), .ZN(n1005) );
  nd02d1 U5982 ( .A1(n6592), .A2(n6361), .ZN(n6376) );
  inv0d0 U5983 ( .I(n11965), .ZN(n2863) );
  inv0d0 U5991 ( .I(n8029), .ZN(n2847) );
  inv0d0 U5992 ( .I(n6137), .ZN(n3563) );
  inv0d0 U5994 ( .I(n9346), .ZN(n3402) );
  nd02d1 U6000 ( .A1(n7453), .A2(n4514), .ZN(n6735) );
  buffd1 U6001 ( .I(n1369), .Z(n1357) );
  nd12d1 U6002 ( .A1(n2615), .A2(n4276), .ZN(n8943) );
  nd02d1 U6005 ( .A1(n8216), .A2(n11373), .ZN(n8965) );
  inv0d0 U6006 ( .I(n5812), .ZN(n4187) );
  inv0d0 U6017 ( .I(n5993), .ZN(n3932) );
  nd02d1 U6021 ( .A1(n6068), .A2(n4692), .ZN(n6077) );
  nd02d1 U6023 ( .A1(n5778), .A2(n8989), .ZN(n8993) );
  inv0d0 U6026 ( .I(n10049), .ZN(n3419) );
  nd02d1 U6029 ( .A1(n4134), .A2(n6652), .ZN(n6819) );
  inv0d1 U6030 ( .I(n1032), .ZN(n1016) );
  inv0d1 U6039 ( .I(n1032), .ZN(n1015) );
  inv0d0 U6040 ( .I(n5084), .ZN(n4029) );
  inv0d1 U6050 ( .I(n1033), .ZN(n1021) );
  inv0d1 U6061 ( .I(n1033), .ZN(n1022) );
  inv0d0 U6062 ( .I(n12038), .ZN(n3510) );
  inv0d0 U6065 ( .I(n9416), .ZN(n3150) );
  nd02d1 U6069 ( .A1(n8050), .A2(n3011), .ZN(n7299) );
  nd02d1 U6072 ( .A1(n4284), .A2(n4330), .ZN(n8968) );
  inv0d0 U6074 ( .I(n6605), .ZN(n3504) );
  nd02d1 U6090 ( .A1(n6058), .A2(n6117), .ZN(n6065) );
  inv0d0 U6092 ( .I(n7327), .ZN(n2830) );
  nd02d1 U6093 ( .A1(n3149), .A2(n5987), .ZN(n11792) );
  inv0d0 U6099 ( .I(n7833), .ZN(n3381) );
  nd12d1 U6101 ( .A1(n24), .A2(n2892), .ZN(n9573) );
  nd04d1 U6108 ( .A1(n1158), .A2(n1443), .A3(n1183), .A4(n1442), .ZN(n24) );
  inv0d0 U6112 ( .I(n7594), .ZN(n4099) );
  inv0d0 U6123 ( .I(n4592), .ZN(n3317) );
  inv0d1 U6126 ( .I(n1031), .ZN(n1028) );
  aoim22d1 U6127 ( .A1(n7935), .A2(n3056), .B1(n11830), .B2(n4729), .Z(n4724)
         );
  inv0d0 U6129 ( .I(n5290), .ZN(n3746) );
  inv0d0 U6130 ( .I(n10707), .ZN(n3744) );
  inv0d0 U6135 ( .I(n11123), .ZN(n2813) );
  inv0d0 U6136 ( .I(n9273), .ZN(n3425) );
  inv0d1 U6138 ( .I(n1034), .ZN(n1024) );
  inv0d1 U6140 ( .I(n1034), .ZN(n1025) );
  nr02d1 U6141 ( .A1(n5521), .A2(n3180), .ZN(n5526) );
  inv0d0 U6142 ( .I(n5528), .ZN(n3180) );
  inv0d1 U6143 ( .I(n1029), .ZN(n999) );
  inv0d0 U6144 ( .I(n4945), .ZN(n4999) );
  inv0d0 U6145 ( .I(n8801), .ZN(n2861) );
  inv0d1 U6146 ( .I(n1034), .ZN(n1026) );
  nd02d1 U6151 ( .A1(n3922), .A2(n3963), .ZN(n6889) );
  inv0d0 U6153 ( .I(n7440), .ZN(n4497) );
  inv0d1 U6158 ( .I(n1034), .ZN(n1027) );
  inv0d0 U6161 ( .I(n9684), .ZN(n4373) );
  inv0d0 U6163 ( .I(n7125), .ZN(n3408) );
  nd02d1 U6164 ( .A1(n3990), .A2(n8870), .ZN(n9099) );
  nd02d1 U6165 ( .A1(n3516), .A2(n5000), .ZN(n8503) );
  inv0d0 U6167 ( .I(n4910), .ZN(n2899) );
  inv0d0 U6169 ( .I(n10941), .ZN(n3301) );
  inv0d1 U6170 ( .I(n1029), .ZN(n1000) );
  nd02d1 U6175 ( .A1(n2837), .A2(n4925), .ZN(n5695) );
  inv0d0 U6176 ( .I(n6583), .ZN(n3213) );
  inv0d0 U6177 ( .I(n6251), .ZN(n3382) );
  inv0d0 U6178 ( .I(n11180), .ZN(n2902) );
  buffd1 U6179 ( .I(n659), .Z(n656) );
  inv0d0 U6181 ( .I(n7132), .ZN(n3406) );
  inv0d0 U6184 ( .I(n7532), .ZN(n4210) );
  nd02d1 U6185 ( .A1(n7454), .A2(n6739), .ZN(n6715) );
  inv0d0 U6187 ( .I(n8766), .ZN(n2995) );
  buffd1 U6191 ( .I(n659), .Z(n657) );
  inv0d0 U6195 ( .I(n5861), .ZN(n4171) );
  nd02d1 U6198 ( .A1(n3514), .A2(n5000), .ZN(n7777) );
  nd02d1 U6199 ( .A1(n6603), .A2(n6204), .ZN(n4535) );
  nd02d1 U6201 ( .A1(n5701), .A2(n5603), .ZN(n5611) );
  inv0d0 U6203 ( .I(n6380), .ZN(n3187) );
  inv0d0 U6207 ( .I(n5379), .ZN(n3477) );
  inv0d0 U6208 ( .I(n8486), .ZN(n3541) );
  buffd1 U6210 ( .I(n1367), .Z(n1362) );
  buffd1 U6211 ( .I(n1367), .Z(n1363) );
  buffd1 U6212 ( .I(n1367), .Z(n1364) );
  inv0d0 U6213 ( .I(n4456), .ZN(n3536) );
  buffd1 U6215 ( .I(n1366), .Z(n1365) );
  buffd1 U6216 ( .I(n1080), .Z(n1059) );
  buffd1 U6217 ( .I(n1369), .Z(n1358) );
  buffd1 U6221 ( .I(n1080), .Z(n1060) );
  buffd1 U6222 ( .I(n1083), .Z(n1051) );
  buffd1 U6223 ( .I(n1081), .Z(n1057) );
  buffd1 U6225 ( .I(n1081), .Z(n1056) );
  inv0d0 U6227 ( .I(n4874), .ZN(n2867) );
  buffd1 U6228 ( .I(n1082), .Z(n1055) );
  buffd1 U6229 ( .I(n1368), .Z(n1361) );
  buffd1 U6230 ( .I(n1369), .Z(n1359) );
  buffd1 U6231 ( .I(n1081), .Z(n1058) );
  buffd1 U6234 ( .I(n1082), .Z(n1054) );
  inv0d0 U6236 ( .I(n4389), .ZN(n4046) );
  buffd1 U6237 ( .I(n1082), .Z(n1053) );
  nd02d1 U6241 ( .A1(n2904), .A2(n2906), .ZN(n10348) );
  buffd1 U6243 ( .I(n1079), .Z(n1062) );
  buffd1 U6246 ( .I(n1078), .Z(n1066) );
  buffd1 U6247 ( .I(n1078), .Z(n1065) );
  buffd1 U6248 ( .I(n1083), .Z(n1052) );
  buffd1 U6249 ( .I(n1368), .Z(n1360) );
  buffd1 U6252 ( .I(n1080), .Z(n1061) );
  buffd1 U6253 ( .I(n1079), .Z(n1064) );
  buffd1 U6258 ( .I(n1079), .Z(n1063) );
  buffd1 U6260 ( .I(n1074), .Z(n1072) );
  buffd1 U6261 ( .I(n1085), .Z(n1044) );
  buffd1 U6263 ( .I(n1077), .Z(n1068) );
  buffd1 U6264 ( .I(n1078), .Z(n1067) );
  inv0d0 U6266 ( .I(n6135), .ZN(n3519) );
  buffd1 U6267 ( .I(n1077), .Z(n1069) );
  buffd1 U6269 ( .I(n1076), .Z(n1070) );
  inv0d0 U6270 ( .I(n5462), .ZN(n3393) );
  buffd1 U6271 ( .I(n1085), .Z(n1045) );
  buffd1 U6272 ( .I(n1085), .Z(n1046) );
  buffd1 U6273 ( .I(n1075), .Z(n1071) );
  buffd1 U6275 ( .I(n1084), .Z(n1047) );
  inv0d0 U6277 ( .I(n5584), .ZN(n3059) );
  buffd1 U6278 ( .I(n1084), .Z(n1048) );
  inv0d0 U6279 ( .I(n9189), .ZN(n3728) );
  buffd1 U6281 ( .I(n1083), .Z(n1050) );
  buffd1 U6282 ( .I(n1084), .Z(n1049) );
  inv0d0 U6283 ( .I(n11373), .ZN(n4260) );
  inv0d0 U6286 ( .I(n4792), .ZN(n2941) );
  inv0d0 U6288 ( .I(n5789), .ZN(n4251) );
  inv0d0 U6292 ( .I(n10138), .ZN(n3184) );
  inv0d0 U6293 ( .I(n4538), .ZN(n3368) );
  inv0d0 U6297 ( .I(n9517), .ZN(n3001) );
  inv0d0 U6301 ( .I(n6549), .ZN(n2844) );
  inv0d0 U6302 ( .I(n7011), .ZN(n3784) );
  inv0d0 U6303 ( .I(n5624), .ZN(n2929) );
  inv0d0 U6305 ( .I(n9363), .ZN(n3388) );
  buffd1 U6306 ( .I(n994), .Z(n992) );
  inv0d0 U6309 ( .I(n9018), .ZN(n4174) );
  buffd1 U6310 ( .I(n996), .Z(n987) );
  buffd1 U6313 ( .I(n996), .Z(n985) );
  buffd1 U6320 ( .I(n995), .Z(n989) );
  buffd1 U6323 ( .I(n995), .Z(n990) );
  buffd1 U6326 ( .I(n996), .Z(n986) );
  buffd1 U6327 ( .I(n994), .Z(n991) );
  inv0d0 U6332 ( .I(n7159), .ZN(n2804) );
  inv0d0 U6334 ( .I(n11543), .ZN(n3937) );
  inv0d0 U6336 ( .I(n8971), .ZN(n4262) );
  buffd1 U6337 ( .I(n995), .Z(n988) );
  inv0d0 U6338 ( .I(n6787), .ZN(n4067) );
  inv0d0 U6339 ( .I(n8132), .ZN(n4835) );
  inv0d0 U6342 ( .I(n12072), .ZN(n4248) );
  inv0d0 U6346 ( .I(n6969), .ZN(n3732) );
  inv0d0 U6348 ( .I(n7316), .ZN(n3003) );
  inv0d0 U6349 ( .I(n6041), .ZN(n2800) );
  inv0d0 U6350 ( .I(n9372), .ZN(n3342) );
  inv0d0 U6351 ( .I(n7884), .ZN(n3191) );
  inv0d0 U6353 ( .I(n8695), .ZN(n3066) );
  inv0d0 U6354 ( .I(n8041), .ZN(n2945) );
  inv0d0 U6356 ( .I(n984), .ZN(n959) );
  inv0d0 U6358 ( .I(n984), .ZN(n960) );
  inv0d0 U6359 ( .I(n4443), .ZN(n3526) );
  inv0d0 U6361 ( .I(n12064), .ZN(n4105) );
  inv0d0 U6362 ( .I(n8850), .ZN(n3377) );
  inv0d0 U6364 ( .I(n7385), .ZN(n3277) );
  inv0d0 U6366 ( .I(n6158), .ZN(n4944) );
  inv0d0 U6369 ( .I(n7769), .ZN(n3514) );
  inv0d0 U6371 ( .I(n6694), .ZN(n5306) );
  inv0d0 U6372 ( .I(n984), .ZN(n961) );
  inv0d0 U6374 ( .I(n5930), .ZN(n4086) );
  inv0d0 U6375 ( .I(n6926), .ZN(n3959) );
  inv0d0 U6377 ( .I(n7736), .ZN(n3779) );
  inv0d0 U6379 ( .I(n5698), .ZN(n5224) );
  inv0d0 U6380 ( .I(n9398), .ZN(n3310) );
  inv0d0 U6383 ( .I(n9354), .ZN(n3379) );
  buffd1 U6385 ( .I(n659), .Z(n658) );
  inv0d0 U6386 ( .I(n7013), .ZN(n3790) );
  inv0d0 U6387 ( .I(n8130), .ZN(n4854) );
  inv0d0 U6388 ( .I(n12016), .ZN(n3412) );
  inv0d0 U6390 ( .I(n10844), .ZN(n3450) );
  inv0d0 U6391 ( .I(n5025), .ZN(n4158) );
  inv0d0 U6392 ( .I(n6944), .ZN(n3890) );
  inv0d0 U6393 ( .I(n6470), .ZN(n3132) );
  inv0d0 U6394 ( .I(n5198), .ZN(n3831) );
  inv0d0 U6397 ( .I(n6711), .ZN(n4272) );
  inv0d0 U6403 ( .I(n11493), .ZN(n4024) );
  inv0d0 U6404 ( .I(n5620), .ZN(n2919) );
  inv0d0 U6405 ( .I(n6128), .ZN(n3529) );
  aoim22d1 U6410 ( .A1(n7866), .A2(n3284), .B1(n8069), .B2(n6320), .Z(n4617)
         );
  buffd1 U6412 ( .I(n1320), .Z(n1319) );
  inv0d0 U6414 ( .I(n7439), .ZN(n4090) );
  inv0d0 U6416 ( .I(n4784), .ZN(n2930) );
  inv0d0 U6418 ( .I(n6815), .ZN(n4101) );
  inv0d0 U6419 ( .I(n12002), .ZN(n3328) );
  inv0d0 U6421 ( .I(n9981), .ZN(n3531) );
  inv0d0 U6423 ( .I(n11367), .ZN(n4229) );
  inv0d0 U6425 ( .I(n7270), .ZN(n3025) );
  inv0d0 U6427 ( .I(n4807), .ZN(n2953) );
  inv0d0 U6429 ( .I(n6217), .ZN(n3373) );
  inv0d0 U6432 ( .I(n7541), .ZN(n4153) );
  inv0d0 U6435 ( .I(n6936), .ZN(n3818) );
  inv0d0 U6437 ( .I(n6686), .ZN(n4230) );
  inv0d0 U6440 ( .I(n8027), .ZN(n2905) );
  inv0d0 U6442 ( .I(n10393), .ZN(n3369) );
  inv0d0 U6443 ( .I(n5424), .ZN(n3360) );
  inv0d0 U6445 ( .I(n8227), .ZN(n4265) );
  inv0d0 U6446 ( .I(n7477), .ZN(n4334) );
  inv0d0 U6447 ( .I(n6647), .ZN(n4735) );
  inv0d0 U6449 ( .I(n7907), .ZN(n3230) );
  inv0d0 U6451 ( .I(n8177), .ZN(n4286) );
  inv0d0 U6455 ( .I(n4458), .ZN(n4441) );
  inv0d0 U6459 ( .I(n8090), .ZN(n3813) );
  inv0d0 U6464 ( .I(n6078), .ZN(n3679) );
  inv0d0 U6468 ( .I(n8973), .ZN(n4283) );
  inv0d0 U6469 ( .I(n5886), .ZN(n4114) );
  inv0d0 U6470 ( .I(n10700), .ZN(n3863) );
  inv0d0 U6471 ( .I(n6378), .ZN(n3178) );
  inv0d0 U6473 ( .I(n7828), .ZN(n3339) );
  inv0d0 U6474 ( .I(n11645), .ZN(n3509) );
  inv0d0 U6476 ( .I(n4897), .ZN(n2839) );
  inv0d0 U6479 ( .I(n9688), .ZN(n4383) );
  inv0d0 U6482 ( .I(n9989), .ZN(n3539) );
  inv0d0 U6484 ( .I(n6492), .ZN(n3101) );
  inv0d0 U6486 ( .I(n10260), .ZN(n2988) );
  inv0d0 U6493 ( .I(n7956), .ZN(n3119) );
  inv0d0 U6498 ( .I(n6781), .ZN(n4065) );
  inv0d0 U6499 ( .I(n9704), .ZN(n4246) );
  inv0d0 U6514 ( .I(n11297), .ZN(n4361) );
  inv0d0 U6518 ( .I(n8848), .ZN(n3400) );
  buffd1 U6530 ( .I(n1172), .Z(n1171) );
  inv0d0 U6534 ( .I(n9626), .ZN(n3806) );
  inv0d0 U6535 ( .I(n5561), .ZN(n3140) );
  inv0d0 U6537 ( .I(n4644), .ZN(n3160) );
  inv0d0 U6538 ( .I(n11362), .ZN(n4270) );
  inv0d0 U6539 ( .I(n6102), .ZN(n3692) );
  inv0d0 U6541 ( .I(n7676), .ZN(n3889) );
  buffd1 U6547 ( .I(n546), .Z(n695) );
  buffd1 U6551 ( .I(n546), .Z(n696) );
  buffd1 U6556 ( .I(n547), .Z(n698) );
  buffd1 U6560 ( .I(n546), .Z(n697) );
  buffd1 U6561 ( .I(n547), .Z(n699) );
  buffd1 U6562 ( .I(n549), .Z(n704) );
  buffd1 U6563 ( .I(n549), .Z(n705) );
  buffd1 U6565 ( .I(n549), .Z(n706) );
  buffd1 U6567 ( .I(n548), .Z(n701) );
  buffd1 U6568 ( .I(n548), .Z(n702) );
  buffd1 U6569 ( .I(n547), .Z(n700) );
  buffd1 U6574 ( .I(n548), .Z(n703) );
  inv0d0 U6577 ( .I(n10051), .ZN(n3333) );
  inv0d0 U6578 ( .I(n11315), .ZN(n4832) );
  buffd1 U6580 ( .I(n1074), .Z(n1073) );
  inv0d0 U6581 ( .I(n8745), .ZN(n3012) );
  inv0d1 U6582 ( .I(n1258), .ZN(n1223) );
  inv0d1 U6583 ( .I(n1258), .ZN(n1224) );
  inv0d0 U6586 ( .I(n8455), .ZN(n3678) );
  inv0d0 U6587 ( .I(n4650), .ZN(n3159) );
  inv0d0 U6588 ( .I(n4490), .ZN(n3502) );
  inv0d0 U6589 ( .I(n8709), .ZN(n2796) );
  inv0d0 U6590 ( .I(n10680), .ZN(n3843) );
  inv0d1 U6591 ( .I(n1031), .ZN(n1006) );
  inv0d0 U6595 ( .I(n6351), .ZN(n3254) );
  inv0d0 U6596 ( .I(n11661), .ZN(n3496) );
  inv0d1 U6598 ( .I(n1031), .ZN(n1007) );
  inv0d1 U6601 ( .I(n1031), .ZN(n1008) );
  inv0d1 U6603 ( .I(n1030), .ZN(n1004) );
  inv0d1 U6604 ( .I(n1030), .ZN(n1002) );
  inv0d1 U6605 ( .I(n1030), .ZN(n1003) );
  inv0d1 U6606 ( .I(n1031), .ZN(n1009) );
  inv0d1 U6608 ( .I(n1031), .ZN(n1010) );
  inv0d0 U6609 ( .I(n7171), .ZN(n3257) );
  inv0d0 U6610 ( .I(n10654), .ZN(n3961) );
  inv0d0 U6611 ( .I(n9700), .ZN(n4243) );
  inv0d0 U6616 ( .I(n8266), .ZN(n4164) );
  inv0d1 U6617 ( .I(n1030), .ZN(n1001) );
  inv0d0 U6618 ( .I(n11909), .ZN(n2835) );
  inv0d0 U6619 ( .I(n5686), .ZN(n2837) );
  inv0d0 U6620 ( .I(n6814), .ZN(n4134) );
  inv0d0 U6621 ( .I(n11784), .ZN(n3149) );
  buffd1 U6622 ( .I(n994), .Z(n993) );
  inv0d1 U6623 ( .I(n1032), .ZN(n1011) );
  inv0d1 U6624 ( .I(n1032), .ZN(n1013) );
  inv0d1 U6625 ( .I(n1032), .ZN(n1012) );
  inv0d1 U6627 ( .I(n1033), .ZN(n1020) );
  inv0d0 U6631 ( .I(n9799), .ZN(n4084) );
  inv0d1 U6633 ( .I(n1032), .ZN(n1014) );
  inv0d0 U6634 ( .I(n6799), .ZN(n4074) );
  inv0d0 U6635 ( .I(n10991), .ZN(n3136) );
  inv0d0 U6638 ( .I(n4410), .ZN(n3792) );
  inv0d0 U6639 ( .I(n7505), .ZN(n4287) );
  inv0d0 U6641 ( .I(n7803), .ZN(n3447) );
  inv0d1 U6642 ( .I(n1033), .ZN(n1019) );
  inv0d1 U6645 ( .I(n1033), .ZN(n1017) );
  inv0d1 U6646 ( .I(n1033), .ZN(n1018) );
  inv0d0 U6649 ( .I(n9758), .ZN(n4223) );
  inv0d0 U6650 ( .I(n8542), .ZN(n3351) );
  inv0d0 U6653 ( .I(n10897), .ZN(n3334) );
  inv0d0 U6654 ( .I(n11797), .ZN(n3148) );
  inv0d0 U6657 ( .I(n7102), .ZN(n3448) );
  inv0d0 U6659 ( .I(n4674), .ZN(n3157) );
  inv0d0 U6660 ( .I(n9279), .ZN(n3493) );
  inv0d0 U6661 ( .I(n9143), .ZN(n3979) );
  inv0d0 U6662 ( .I(n6020), .ZN(n3829) );
  inv0d0 U6663 ( .I(n10450), .ZN(n4580) );
  inv0d0 U6664 ( .I(n11257), .ZN(n3860) );
  inv0d0 U6666 ( .I(n8718), .ZN(n3083) );
  inv0d0 U6667 ( .I(n5151), .ZN(n3931) );
  inv0d0 U6668 ( .I(n11221), .ZN(n3135) );
  inv0d0 U6669 ( .I(n8465), .ZN(n3525) );
  inv0d0 U6670 ( .I(n8930), .ZN(n4227) );
  inv0d0 U6677 ( .I(n5940), .ZN(n4087) );
  inv0d1 U6683 ( .I(n1029), .ZN(n998) );
  inv0d1 U6688 ( .I(n1034), .ZN(n1023) );
  inv0d0 U6689 ( .I(n7364), .ZN(n3067) );
  inv0d0 U6690 ( .I(n8669), .ZN(n3018) );
  inv0d0 U6694 ( .I(n10883), .ZN(n3376) );
  inv0d0 U6697 ( .I(n4937), .ZN(n2987) );
  inv0d0 U6698 ( .I(n7598), .ZN(n4094) );
  inv0d0 U6702 ( .I(n9555), .ZN(n2857) );
  inv0d0 U6703 ( .I(n6210), .ZN(n3415) );
  inv0d0 U6704 ( .I(n7137), .ZN(n3380) );
  inv0d0 U6708 ( .I(n7486), .ZN(n4366) );
  nr02d1 U6710 ( .A1(n3685), .A2(N5285), .ZN(n3651) );
  nd02d1 U6718 ( .A1(N3884), .A2(n949), .ZN(n3609) );
  nd02d1 U6719 ( .A1(n4237), .A2(n4254), .ZN(n4242) );
  inv0d0 U6720 ( .I(n4240), .ZN(n2757) );
  buffd1 U6729 ( .I(n4245), .Z(n496) );
  nd03d1 U6730 ( .A1(n4242), .A2(n2778), .A3(n4235), .ZN(n4245) );
  oai211d1 U6731 ( .C1(n3655), .C2(n3689), .A(n493), .B(n2771), .ZN(n3677) );
  inv0d0 U6733 ( .I(n499), .ZN(n500) );
  inv0d0 U6745 ( .I(n501), .ZN(n502) );
  inv0d0 U6746 ( .I(n503), .ZN(n504) );
  inv0d0 U6747 ( .I(n505), .ZN(n506) );
  inv0d0 U6754 ( .I(n507), .ZN(n508) );
  inv0d0 U6755 ( .I(n418), .ZN(n509) );
  inv0d0 U6756 ( .I(n419), .ZN(n510) );
  inv0d0 U6757 ( .I(n512), .ZN(n513) );
  inv0d0 U6758 ( .I(n3687), .ZN(n2755) );
  nr02d1 U6759 ( .A1(n3685), .A2(n3655), .ZN(n3688) );
  inv0d0 U6761 ( .I(n3657), .ZN(n2771) );
  inv0d0 U6762 ( .I(n2730), .ZN(n2743) );
  nd03d1 U6765 ( .A1(n3825), .A2(n12206), .A3(n3794), .ZN(n3797) );
  nr02d1 U6768 ( .A1(n3657), .A2(n4254), .ZN(n3707) );
  nd03d1 U6772 ( .A1(n3825), .A2(n2786), .A3(n3794), .ZN(n3710) );
  nd03d1 U6776 ( .A1(n3825), .A2(n2786), .A3(n4010), .ZN(n3980) );
  nd03d1 U6777 ( .A1(n3884), .A2(n2785), .A3(n4010), .ZN(n4100) );
  nd03d1 U6779 ( .A1(n3796), .A2(n12206), .A3(n4010), .ZN(n4069) );
  nd03d1 U6780 ( .A1(n3884), .A2(n12207), .A3(n4010), .ZN(n4131) );
  nd03d1 U6781 ( .A1(n3948), .A2(n12207), .A3(n4010), .ZN(n4194) );
  nd03d1 U6784 ( .A1(n3825), .A2(n12206), .A3(n4010), .ZN(n4040) );
  nd03d1 U6785 ( .A1(n3796), .A2(n2786), .A3(n4010), .ZN(n4011) );
  nd03d1 U6795 ( .A1(n3948), .A2(n2785), .A3(n4010), .ZN(n4162) );
  nd03d1 U6796 ( .A1(n2775), .A2(n2779), .A3(n495), .ZN(n3662) );
  nd02d1 U6797 ( .A1(n2759), .A2(n3682), .ZN(n3658) );
  inv0d0 U6798 ( .I(n511), .ZN(N4664) );
  nd03d1 U6804 ( .A1(n3794), .A2(n2785), .A3(n3948), .ZN(n3918) );
  nd03d1 U6805 ( .A1(n3794), .A2(n12207), .A3(n3884), .ZN(n3885) );
  nd03d1 U6806 ( .A1(n3794), .A2(n2786), .A3(n3796), .ZN(n3767) );
  nd03d1 U6807 ( .A1(n3794), .A2(n2785), .A3(n3884), .ZN(n3855) );
  nd03d1 U6813 ( .A1(n3794), .A2(n12207), .A3(n3948), .ZN(n3949) );
  nd03d1 U6822 ( .A1(n3794), .A2(n12206), .A3(n3796), .ZN(n3827) );
  inv0d2 U6825 ( .I(n956), .ZN(n955) );
  buffd1 U6826 ( .I(n4363), .Z(n754) );
  buffd1 U6827 ( .I(n4367), .Z(n738) );
  buffd1 U6830 ( .I(n4359), .Z(n773) );
  buffd1 U6831 ( .I(n4360), .Z(n767) );
  buffd1 U6833 ( .I(n4372), .Z(n712) );
  buffd1 U6836 ( .I(n4370), .Z(n725) );
  buffd1 U6837 ( .I(n4356), .Z(n797) );
  buffd1 U6840 ( .I(n4353), .Z(n810) );
  buffd1 U6841 ( .I(n739), .Z(n743) );
  buffd1 U6842 ( .I(n4367), .Z(n739) );
  buffd1 U6844 ( .I(n755), .Z(n759) );
  buffd1 U6846 ( .I(n4363), .Z(n755) );
  buffd1 U6849 ( .I(n713), .Z(n717) );
  buffd1 U6864 ( .I(n4372), .Z(n713) );
  buffd1 U6868 ( .I(n811), .Z(n815) );
  buffd1 U6871 ( .I(n4353), .Z(n811) );
  buffd1 U6877 ( .I(n774), .Z(n778) );
  buffd1 U6878 ( .I(n4359), .Z(n774) );
  buffd1 U6879 ( .I(n768), .Z(n772) );
  buffd1 U6880 ( .I(n4360), .Z(n768) );
  buffd1 U6885 ( .I(n726), .Z(n730) );
  buffd1 U6888 ( .I(n4370), .Z(n726) );
  buffd1 U6890 ( .I(n798), .Z(n802) );
  buffd1 U6891 ( .I(n4356), .Z(n798) );
  nd02d1 U6893 ( .A1(n4337), .A2(n495), .ZN(n4335) );
  buffd1 U6894 ( .I(n3680), .Z(n495) );
  nr02d1 U6899 ( .A1(n3667), .A2(n3654), .ZN(n3680) );
  nd02d1 U6900 ( .A1(n4329), .A2(n495), .ZN(n4327) );
  nd02d1 U6902 ( .A1(n4337), .A2(n2), .ZN(n4364) );
  buffd1 U6903 ( .I(n2765), .Z(n538) );
  buffd1 U6904 ( .I(n2765), .Z(n539) );
  buffd1 U6911 ( .I(n2765), .Z(n540) );
  buffd1 U6912 ( .I(n2760), .Z(n542) );
  buffd1 U6917 ( .I(n2760), .Z(n543) );
  buffd1 U6923 ( .I(n2760), .Z(n544) );
  buffd1 U6926 ( .I(n2763), .Z(n526) );
  buffd1 U6927 ( .I(n2763), .Z(n527) );
  buffd1 U6929 ( .I(n2763), .Z(n528) );
  buffd1 U6932 ( .I(n2764), .Z(n530) );
  buffd1 U6936 ( .I(n2764), .Z(n531) );
  buffd1 U6941 ( .I(n2764), .Z(n532) );
  buffd1 U6945 ( .I(n2765), .Z(n534) );
  buffd1 U6947 ( .I(n2765), .Z(n535) );
  buffd1 U6955 ( .I(n2765), .Z(n536) );
  buffd1 U6958 ( .I(n2761), .Z(n518) );
  buffd1 U6965 ( .I(n2761), .Z(n519) );
  buffd1 U6972 ( .I(n2761), .Z(n520) );
  buffd1 U6974 ( .I(n2762), .Z(n522) );
  buffd1 U6981 ( .I(n2762), .Z(n523) );
  buffd1 U6994 ( .I(n2762), .Z(n524) );
  buffd1 U6995 ( .I(n2760), .Z(n514) );
  buffd1 U6996 ( .I(n2760), .Z(n515) );
  buffd1 U7002 ( .I(n2760), .Z(n516) );
  buffd1 U7004 ( .I(n537), .Z(n541) );
  buffd1 U7005 ( .I(n517), .Z(n545) );
  buffd1 U7006 ( .I(n2763), .Z(n529) );
  buffd1 U7009 ( .I(n2764), .Z(n533) );
  buffd1 U7010 ( .I(n2765), .Z(n537) );
  buffd1 U7011 ( .I(n2761), .Z(n521) );
  buffd1 U7012 ( .I(n2762), .Z(n525) );
  buffd1 U7013 ( .I(n2760), .Z(n517) );
  nd02d1 U7014 ( .A1(n4329), .A2(n2), .ZN(n4358) );
  inv0d0 U7017 ( .I(n3588), .ZN(n2777) );
  nd02d1 U7019 ( .A1(n497), .A2(N26489), .ZN(n3706) );
  nr02d1 U7020 ( .A1(n3656), .A2(N3855), .ZN(n3652) );
  inv0d0 U7023 ( .I(N26489), .ZN(n2783) );
  nr02d1 U7025 ( .A1(n3646), .A2(n3588), .ZN(n3589) );
  inv0d0 U7027 ( .I(n1411), .ZN(n1420) );
  inv0d0 U7029 ( .I(N26480), .ZN(n2781) );
  nd02d1 U7032 ( .A1(n4206), .A2(n4197), .ZN(n3716) );
  nd02d1 U7033 ( .A1(n4193), .A2(n4197), .ZN(n3720) );
  nd02d1 U7034 ( .A1(n4208), .A2(n4197), .ZN(n3718) );
  nd02d1 U7036 ( .A1(n4204), .A2(n4197), .ZN(n3714) );
  nd02d1 U7037 ( .A1(n4200), .A2(n4197), .ZN(n3711) );
  nd02d1 U7039 ( .A1(n4202), .A2(n4197), .ZN(n3713) );
  nd02d1 U7040 ( .A1(n4192), .A2(n4198), .ZN(n3754) );
  nd02d1 U7041 ( .A1(n4221), .A2(n4198), .ZN(n3739) );
  nd02d1 U7042 ( .A1(n4212), .A2(n4198), .ZN(n3724) );
  nd02d1 U7044 ( .A1(n4221), .A2(n4206), .ZN(n3747) );
  nd02d1 U7051 ( .A1(n4212), .A2(n4206), .ZN(n3731) );
  nd02d1 U7052 ( .A1(n4192), .A2(n4202), .ZN(n3758) );
  nd02d1 U7053 ( .A1(n4221), .A2(n4202), .ZN(n3743) );
  nd02d1 U7057 ( .A1(n4212), .A2(n4202), .ZN(n3727) );
  nd02d1 U7060 ( .A1(n4192), .A2(n4208), .ZN(n3763) );
  nd02d1 U7061 ( .A1(n4212), .A2(n4208), .ZN(n3733) );
  nd02d1 U7063 ( .A1(n4221), .A2(n4193), .ZN(n3750) );
  nd02d1 U7065 ( .A1(n4212), .A2(n4193), .ZN(n3735) );
  nd02d1 U7066 ( .A1(n4192), .A2(n4193), .ZN(n3765) );
  nd02d1 U7071 ( .A1(n4192), .A2(n4204), .ZN(n3760) );
  nd02d1 U7074 ( .A1(n4221), .A2(n4204), .ZN(n3745) );
  nd02d1 U7076 ( .A1(n4212), .A2(n4204), .ZN(n3729) );
  nd02d1 U7080 ( .A1(n4192), .A2(n4200), .ZN(n3756) );
  nd02d1 U7082 ( .A1(n4221), .A2(n4200), .ZN(n3741) );
  nd02d1 U7083 ( .A1(n4197), .A2(n4198), .ZN(n3709) );
  nd02d1 U7084 ( .A1(n4192), .A2(n4206), .ZN(n3762) );
  nd02d1 U7086 ( .A1(n4221), .A2(n4208), .ZN(n3749) );
  nd02d1 U7087 ( .A1(n4211), .A2(n4197), .ZN(n3768) );
  nd02d1 U7090 ( .A1(n4211), .A2(n4212), .ZN(n3722) );
  nd02d1 U7096 ( .A1(n4212), .A2(n4200), .ZN(n3726) );
  nd02d1 U7099 ( .A1(n4192), .A2(n4211), .ZN(n3752) );
  nd02d1 U7100 ( .A1(n4221), .A2(n4211), .ZN(n3737) );
  inv0d0 U7101 ( .I(N29414), .ZN(N3212) );
  nr02d1 U7102 ( .A1(n3654), .A2(N3855), .ZN(n3646) );
  nd02d1 U7104 ( .A1(n2781), .A2(n2776), .ZN(n3670) );
  inv0d0 U7110 ( .I(n9175), .ZN(n3871) );
  nd03d1 U7111 ( .A1(n6681), .A2(n4376), .A3(n4384), .ZN(n6672) );
  inv0d0 U7114 ( .I(n9497), .ZN(n2936) );
  nr02d1 U7117 ( .A1(n5959), .A2(n8204), .ZN(n6719) );
  nr02d1 U7118 ( .A1(n3129), .A2(n7258), .ZN(n6430) );
  nr02d1 U7123 ( .A1(n5420), .A2(n10847), .ZN(n6194) );
  nr02d1 U7124 ( .A1(n6174), .A2(n3577), .ZN(n5345) );
  inv0d0 U7127 ( .I(n10671), .ZN(n3815) );
  inv0d0 U7130 ( .I(n10334), .ZN(n2823) );
  inv0d0 U7133 ( .I(n4641), .ZN(n3170) );
  nr02d1 U7134 ( .A1(n6589), .A2(n12072), .ZN(n8197) );
  nd02d1 U7135 ( .A1(n7319), .A2(n5126), .ZN(n11866) );
  nr02d1 U7136 ( .A1(n6948), .A2(n5775), .ZN(n5890) );
  inv0d0 U7137 ( .I(n4548), .ZN(n3370) );
  nr02d1 U7138 ( .A1(n4554), .A2(n11705), .ZN(n11704) );
  inv0d0 U7140 ( .I(n9136), .ZN(n3978) );
  inv0d0 U7141 ( .I(n8792), .ZN(n2817) );
  nr02d1 U7142 ( .A1(n6747), .A2(n5527), .ZN(n4985) );
  nr02d1 U7144 ( .A1(n7985), .A2(n2985), .ZN(n10257) );
  inv0d0 U7146 ( .I(n11970), .ZN(n2985) );
  nd02d1 U7147 ( .A1(n3402), .A2(n3375), .ZN(n12008) );
  inv0d0 U7150 ( .I(n1842), .ZN(N12898) );
  inv0d0 U7151 ( .I(n1841), .ZN(n1843) );
  nd02d1 U7153 ( .A1(n4821), .A2(n4820), .ZN(n11876) );
  nr02d1 U7155 ( .A1(n5034), .A2(n9436), .ZN(n11220) );
  nr02d1 U7156 ( .A1(n7019), .A2(n10697), .ZN(n11256) );
  nr02d1 U7157 ( .A1(n10773), .A2(n7028), .ZN(n5745) );
  nr02d1 U7158 ( .A1(n6993), .A2(n5806), .ZN(n4960) );
  nr02d1 U7159 ( .A1(n6481), .A2(n6930), .ZN(n12059) );
  nr02d1 U7161 ( .A1(n5221), .A2(n10282), .ZN(n10288) );
  nr02d1 U7164 ( .A1(n6291), .A2(n7882), .ZN(n7227) );
  nr02d1 U7167 ( .A1(n3577), .A2(n7015), .ZN(n11622) );
  nr02d1 U7170 ( .A1(n7428), .A2(n6917), .ZN(n6003) );
  nr02d1 U7171 ( .A1(n6550), .A2(n5110), .ZN(n7455) );
  nr02d1 U7173 ( .A1(n6538), .A2(n5063), .ZN(n7003) );
  nr02d1 U7174 ( .A1(n7319), .A2(n7316), .ZN(n4814) );
  nr02d1 U7176 ( .A1(n9606), .A2(n6346), .ZN(n4972) );
  nr02d1 U7177 ( .A1(n4979), .A2(n7222), .ZN(n5720) );
  nr02d1 U7179 ( .A1(n11378), .A2(n8222), .ZN(n8988) );
  nr02d1 U7180 ( .A1(n6400), .A2(n4745), .ZN(n6657) );
  inv0d0 U7181 ( .I(n1754), .ZN(n1756) );
  nr02d1 U7183 ( .A1(n7155), .A2(n6038), .ZN(n7685) );
  nr02d1 U7185 ( .A1(n6297), .A2(n4427), .ZN(n6602) );
  nr02d1 U7189 ( .A1(n4), .A2(n8563), .ZN(n6232) );
  nr02d1 U7191 ( .A1(n10405), .A2(n6923), .ZN(n4442) );
  nr02d1 U7194 ( .A1(n6207), .A2(n4292), .ZN(n8126) );
  nr02d1 U7197 ( .A1(n11561), .A2(n6016), .ZN(n6013) );
  nr02d1 U7199 ( .A1(n5897), .A2(n9050), .ZN(n6787) );
  nr02d1 U7201 ( .A1(n4119), .A2(n5876), .ZN(n11430) );
  nr02d1 U7203 ( .A1(n5504), .A2(n11770), .ZN(n10106) );
  inv0d0 U7205 ( .I(n11026), .ZN(n2812) );
  nd02d1 U7206 ( .A1(n8798), .A2(n5604), .ZN(n10297) );
  nr02d1 U7208 ( .A1(n10413), .A2(n6938), .ZN(n5780) );
  inv0d0 U7213 ( .I(n7206), .ZN(n3256) );
  nr02d1 U7215 ( .A1(n6160), .A2(n3129), .ZN(n5706) );
  nr02d1 U7220 ( .A1(n7690), .A2(n11259), .ZN(n5219) );
  aoim22d1 U7221 ( .A1(n3529), .A2(n4445), .B1(n4446), .B2(n4442), .Z(n4440)
         );
  nr02d1 U7222 ( .A1(n5004), .A2(n5005), .ZN(n4447) );
  nr02d1 U7223 ( .A1(n8766), .A2(n9525), .ZN(n11972) );
  nr02d1 U7224 ( .A1(n6586), .A2(n5204), .ZN(n6663) );
  nr02d1 U7225 ( .A1(n6548), .A2(n5106), .ZN(n5852) );
  inv0d0 U7226 ( .I(n5847), .ZN(n4506) );
  nr02d1 U7227 ( .A1(n6246), .A2(n4313), .ZN(n8857) );
  nr02d1 U7231 ( .A1(n6330), .A2(n4491), .ZN(n5077) );
  nr02d1 U7232 ( .A1(n4671), .A2(n11984), .ZN(n5529) );
  nr02d1 U7233 ( .A1(n6119), .A2(n6935), .ZN(n5767) );
  nr02d1 U7234 ( .A1(n6024), .A2(n6388), .ZN(n6134) );
  nr02d1 U7235 ( .A1(n12068), .A2(n10537), .ZN(n7548) );
  nd02d1 U7236 ( .A1(n3399), .A2(n5046), .ZN(n12006) );
  nr02d1 U7238 ( .A1(n6445), .A2(n8572), .ZN(n5463) );
  inv0d0 U7242 ( .I(n6283), .ZN(n3329) );
  inv0d0 U7244 ( .I(n7161), .ZN(n3325) );
  inv0d0 U7246 ( .I(n7950), .ZN(n3068) );
  inv0d0 U7247 ( .I(n8259), .ZN(n4159) );
  nr02d1 U7250 ( .A1(n8082), .A2(n7711), .ZN(n5271) );
  nr02d1 U7251 ( .A1(n11186), .A2(n11187), .ZN(n9563) );
  nr02d1 U7256 ( .A1(n7047), .A2(n11330), .ZN(n11333) );
  inv0d0 U7257 ( .I(n1687), .ZN(n1688) );
  nr02d1 U7262 ( .A1(n9227), .A2(n10746), .ZN(n5331) );
  nr02d1 U7266 ( .A1(n6593), .A2(n6594), .ZN(n6350) );
  inv0d0 U7267 ( .I(n5070), .ZN(n4021) );
  nr02d1 U7268 ( .A1(n7182), .A2(n6748), .ZN(n6665) );
  nr02d1 U7269 ( .A1(n6707), .A2(n5466), .ZN(n7487) );
  nr02d1 U7270 ( .A1(n7183), .A2(n6070), .ZN(n6702) );
  nd03d1 U7271 ( .A1(n3114), .A2(n9601), .A3(n3081), .ZN(n9476) );
  inv0d0 U7274 ( .I(n4546), .ZN(n3349) );
  nr02d1 U7277 ( .A1(n8096), .A2(n5851), .ZN(n5783) );
  nr02d1 U7279 ( .A1(n7022), .A2(n11552), .ZN(n10657) );
  inv0d0 U7282 ( .I(n5210), .ZN(n3842) );
  inv0d0 U7283 ( .I(n5921), .ZN(n4107) );
  inv0d0 U7284 ( .I(n11935), .ZN(n2833) );
  inv0d0 U7285 ( .I(n11620), .ZN(n2791) );
  nd02d1 U7289 ( .A1(n3684), .A2(n5345), .ZN(n6125) );
  inv0d0 U7290 ( .I(n8362), .ZN(n2794) );
  inv0d0 U7294 ( .I(n6740), .ZN(n4328) );
  nr02d1 U7295 ( .A1(n11716), .A2(n8850), .ZN(n4559) );
  nr02d1 U7297 ( .A1(n4394), .A2(n4433), .ZN(n5170) );
  nr02d1 U7299 ( .A1(n5106), .A2(n4174), .ZN(n11416) );
  nr02d1 U7300 ( .A1(n6750), .A2(n5816), .ZN(n5821) );
  nr02d1 U7301 ( .A1(n11182), .A2(n10343), .ZN(n4910) );
  inv0d0 U7302 ( .I(n4525), .ZN(n3361) );
  nr02d1 U7305 ( .A1(n6411), .A2(n4754), .ZN(n6697) );
  nr02d1 U7306 ( .A1(n8704), .A2(n6287), .ZN(n11833) );
  aoim22d1 U7307 ( .A1(n3956), .A2(n3814), .B1(n9892), .B2(n3821), .Z(n12061)
         );
  inv0d0 U7309 ( .I(N9484), .ZN(n7603) );
  inv0d0 U7312 ( .I(n8988), .ZN(n4267) );
  inv0d0 U7315 ( .I(n5304), .ZN(n3700) );
  nr02d1 U7316 ( .A1(n5631), .A2(n6296), .ZN(n4977) );
  nr02d1 U7318 ( .A1(n8208), .A2(n11368), .ZN(n7511) );
  inv0d0 U7321 ( .I(n8264), .ZN(n4218) );
  nr02d1 U7322 ( .A1(n6823), .A2(n6825), .ZN(n9081) );
  inv0d0 U7324 ( .I(n11324), .ZN(n4575) );
  nr02d1 U7325 ( .A1(n11877), .A2(n10258), .ZN(n4826) );
  inv0d0 U7326 ( .I(n6681), .ZN(n4551) );
  inv0d0 U7327 ( .I(n11705), .ZN(n3346) );
  inv0d0 U7328 ( .I(n4547), .ZN(n3371) );
  nr02d1 U7329 ( .A1(n6146), .A2(n10472), .ZN(n11338) );
  nr02d1 U7332 ( .A1(n6056), .A2(n5899), .ZN(n8282) );
  nr02d1 U7334 ( .A1(n7121), .A2(n11828), .ZN(n8691) );
  nr02d1 U7336 ( .A1(n6896), .A2(n5144), .ZN(n8356) );
  nr02d1 U7337 ( .A1(n6229), .A2(n5504), .ZN(n6333) );
  inv0d0 U7338 ( .I(n6546), .ZN(n2843) );
  nd03d1 U7343 ( .A1(n3542), .A2(n3558), .A3(n6141), .ZN(n6136) );
  aoim22d1 U7345 ( .A1(n6148), .A2(n6149), .B1(n6150), .B2(n5363), .Z(n6142)
         );
  nd02d1 U7346 ( .A1(n7315), .A2(n5607), .ZN(n11864) );
  inv0d0 U7348 ( .I(n6431), .ZN(n3226) );
  nr02d1 U7350 ( .A1(n6469), .A2(n9622), .ZN(n9232) );
  inv0d0 U7356 ( .I(n11757), .ZN(n3264) );
  inv0d0 U7358 ( .I(n5628), .ZN(n2923) );
  nr02d1 U7360 ( .A1(n8658), .A2(n6588), .ZN(n6583) );
  nr02d1 U7362 ( .A1(n6143), .A2(n9259), .ZN(n9255) );
  inv0d0 U7363 ( .I(n10039), .ZN(n3441) );
  inv0d0 U7366 ( .I(n5273), .ZN(n3699) );
  inv0d0 U7367 ( .I(n8508), .ZN(n3497) );
  inv0d0 U7369 ( .I(n8520), .ZN(n3498) );
  inv0d0 U7370 ( .I(n6188), .ZN(n3420) );
  nd02d1 U7372 ( .A1(n11993), .A2(n5515), .ZN(n11785) );
  inv0d0 U7374 ( .I(n6893), .ZN(n3923) );
  inv0d0 U7376 ( .I(n9078), .ZN(n4136) );
  inv0d0 U7377 ( .I(n8176), .ZN(n4226) );
  inv0d0 U7379 ( .I(n5781), .ZN(n3912) );
  inv0d0 U7382 ( .I(n11061), .ZN(n3019) );
  nr02d1 U7384 ( .A1(n5146), .A2(n11746), .ZN(n11751) );
  nd03d1 U7385 ( .A1(n5219), .A2(n9909), .A3(n3840), .ZN(n9908) );
  inv0d0 U7388 ( .I(n9914), .ZN(n3811) );
  nd03d1 U7389 ( .A1(n6494), .A2(n6500), .A3(n6501), .ZN(n6498) );
  nr02d1 U7391 ( .A1(n4993), .A2(n10045), .ZN(n9319) );
  inv0d0 U7394 ( .I(n4919), .ZN(n5482) );
  nr02d1 U7395 ( .A1(n5046), .A2(n11716), .ZN(n6247) );
  inv0d0 U7397 ( .I(n4812), .ZN(n3000) );
  inv0d0 U7398 ( .I(n7626), .ZN(n4030) );
  nr02d1 U7399 ( .A1(n7245), .A2(n8311), .ZN(n11473) );
  inv0d0 U7400 ( .I(n7515), .ZN(n4288) );
  inv0d0 U7403 ( .I(n10553), .ZN(n4120) );
  inv0d0 U7406 ( .I(n7812), .ZN(n3422) );
  nr02d1 U7407 ( .A1(n5839), .A2(n6250), .ZN(n8862) );
  nr02d1 U7411 ( .A1(n5193), .A2(n11556), .ZN(n6936) );
  inv0d0 U7413 ( .I(n4705), .ZN(n3033) );
  nr02d1 U7414 ( .A1(n8813), .A2(n4919), .ZN(n11937) );
  nr02d1 U7417 ( .A1(n6646), .A2(n5312), .ZN(n8119) );
  nd02d1 U7418 ( .A1(n5718), .A2(n5719), .ZN(n5502) );
  nr02d1 U7420 ( .A1(n6240), .A2(n9304), .ZN(n10837) );
  nr02d1 U7422 ( .A1(n5371), .A2(n6151), .ZN(n6154) );
  nr02d1 U7425 ( .A1(n8873), .A2(n5936), .ZN(n6652) );
  inv0d0 U7427 ( .I(n8052), .ZN(n3091) );
  nr02d1 U7432 ( .A1(n6268), .A2(n4326), .ZN(n6661) );
  inv0d0 U7433 ( .I(n5761), .ZN(n3849) );
  nr02d1 U7434 ( .A1(n6428), .A2(n11062), .ZN(n11854) );
  inv0d0 U7435 ( .I(n9232), .ZN(n3715) );
  nd03d1 U7439 ( .A1(n9232), .A2(n5345), .A3(n9236), .ZN(n9233) );
  nd02d1 U7440 ( .A1(N10836), .A2(n6955), .ZN(n5227) );
  nr02d1 U7442 ( .A1(n6200), .A2(n4222), .ZN(n8884) );
  nr02d1 U7443 ( .A1(n6667), .A2(n5831), .ZN(n5042) );
  nr02d1 U7444 ( .A1(n6198), .A2(n10850), .ZN(n5424) );
  inv0d0 U7446 ( .I(n10657), .ZN(n3954) );
  inv0d0 U7449 ( .I(n7861), .ZN(n2799) );
  nr02d1 U7451 ( .A1(n5775), .A2(n7572), .ZN(n5888) );
  inv0d0 U7453 ( .I(n9311), .ZN(n3492) );
  nr02d1 U7454 ( .A1(n9638), .A2(n11277), .ZN(n6648) );
  nd02d1 U7456 ( .A1(n9563), .A2(n10312), .ZN(n10311) );
  nr02d1 U7457 ( .A1(n6894), .A2(n5727), .ZN(n8039) );
  nd02d1 U7458 ( .A1(n8670), .A2(n6437), .ZN(n7258) );
  nd03d1 U7459 ( .A1(n11103), .A2(n6512), .A3(n9526), .ZN(n11106) );
  inv0d0 U7460 ( .I(n4708), .ZN(n3039) );
  nr02d1 U7461 ( .A1(n8208), .A2(n4253), .ZN(n6721) );
  nr02d1 U7462 ( .A1(n6654), .A2(n5320), .ZN(n4914) );
  nr02d1 U7463 ( .A1(n6077), .A2(n5296), .ZN(n6078) );
  nr02d1 U7464 ( .A1(n5766), .A2(n5276), .ZN(n7422) );
  nr02d1 U7465 ( .A1(n8863), .A2(n5234), .ZN(n5759) );
  nr02d1 U7467 ( .A1(n10952), .A2(n5500), .ZN(n6331) );
  nr02d1 U7471 ( .A1(n7121), .A2(n5980), .ZN(n4730) );
  nr02d1 U7473 ( .A1(n11857), .A2(n9504), .ZN(n4792) );
  nr02d1 U7474 ( .A1(n6519), .A2(n5003), .ZN(n4945) );
  or02d0 U7479 ( .A1(n7215), .A2(n1727), .Z(n6364) );
  nr02d1 U7480 ( .A1(n5957), .A2(n7442), .ZN(n7440) );
  nr02d1 U7481 ( .A1(n7413), .A2(n8858), .ZN(n5752) );
  nr02d1 U7483 ( .A1(n5153), .A2(n7430), .ZN(n6902) );
  nr02d1 U7485 ( .A1(n4871), .A2(n6653), .ZN(n8897) );
  nr02d1 U7487 ( .A1(n6778), .A2(n5573), .ZN(n5082) );
  nd12d1 U7489 ( .A1(n11156), .A2(n2885), .ZN(n4920) );
  nr02d1 U7490 ( .A1(n7599), .A2(n6830), .ZN(n5024) );
  nr02d1 U7491 ( .A1(n5558), .A2(n5167), .ZN(n6910) );
  nr02d1 U7492 ( .A1(n6305), .A2(n4450), .ZN(n9246) );
  nr02d1 U7493 ( .A1(n5757), .A2(n5256), .ZN(n11583) );
  nr02d1 U7494 ( .A1(n9714), .A2(n6713), .ZN(n5789) );
  nr02d1 U7496 ( .A1(n6990), .A2(n5802), .ZN(n6561) );
  nr02d1 U7497 ( .A1(n7069), .A2(n5927), .ZN(n5724) );
  nr02d1 U7502 ( .A1(n9982), .A2(n12042), .ZN(n9977) );
  nd02d1 U7504 ( .A1(N13570), .A2(n10958), .ZN(n6593) );
  nr02d1 U7505 ( .A1(n5146), .A2(n5485), .ZN(n11752) );
  nr02d1 U7506 ( .A1(n6508), .A2(n4980), .ZN(n4917) );
  nd12d1 U7508 ( .A1(n25), .A2(n4804), .ZN(n7316) );
  nd04d1 U7512 ( .A1(n1342), .A2(n1299), .A3(n1246), .A4(n1541), .ZN(n25) );
  nr02d1 U7513 ( .A1(n5322), .A2(n6982), .ZN(n9539) );
  nr02d1 U7514 ( .A1(n6670), .A2(n5397), .ZN(n7388) );
  nr02d1 U7515 ( .A1(n6613), .A2(n6172), .ZN(n5384) );
  nr02d1 U7517 ( .A1(n5728), .A2(n7918), .ZN(n8680) );
  nr02d1 U7518 ( .A1(n7176), .A2(n6056), .ZN(n6656) );
  nr02d1 U7521 ( .A1(n11619), .A2(n7411), .ZN(n8453) );
  nr02d1 U7523 ( .A1(n7104), .A2(n5958), .ZN(n7450) );
  nr02d1 U7524 ( .A1(n5242), .A2(n3246), .ZN(n10969) );
  nr02d1 U7528 ( .A1(n6507), .A2(n9688), .ZN(n11336) );
  nr02d1 U7530 ( .A1(n5109), .A2(n7645), .ZN(n7648) );
  nr02d1 U7532 ( .A1(n3907), .A2(n9119), .ZN(n9121) );
  inv0d0 U7534 ( .I(n5953), .ZN(n3984) );
  nr02d1 U7538 ( .A1(n9573), .A2(n9574), .ZN(n4898) );
  nr02d1 U7542 ( .A1(n8093), .A2(n5139), .ZN(n8092) );
  nr02d1 U7543 ( .A1(n5251), .A2(n5757), .ZN(n5261) );
  nr02d1 U7544 ( .A1(n6825), .A2(n7034), .ZN(n6651) );
  nd02d1 U7546 ( .A1(N14882), .A2(n8763), .ZN(n8766) );
  nr02d1 U7547 ( .A1(n7075), .A2(n5933), .ZN(n5002) );
  nr02d1 U7550 ( .A1(n6254), .A2(n6253), .ZN(n6251) );
  inv0d0 U7551 ( .I(n8844), .ZN(n3162) );
  inv0d0 U7553 ( .I(n8604), .ZN(n3258) );
  inv0d0 U7554 ( .I(n6057), .ZN(n3859) );
  nd02d1 U7556 ( .A1(N13778), .A2(n11992), .ZN(n6379) );
  aoim22d1 U7557 ( .A1(n4031), .A2(n6862), .B1(n6863), .B2(n4389), .Z(n6859)
         );
  inv0d0 U7558 ( .I(n7437), .ZN(n4031) );
  aoim22d1 U7561 ( .A1(n6299), .A2(n6300), .B1(n6301), .B2(n6302), .Z(n6288)
         );
  inv0d0 U7562 ( .I(n6292), .ZN(n3324) );
  nd03d1 U7563 ( .A1(n5744), .A2(n5745), .A3(n3523), .ZN(n5352) );
  nr02d1 U7564 ( .A1(n7774), .A2(n6100), .ZN(n5000) );
  nd02d1 U7567 ( .A1(n3369), .A2(n10065), .ZN(n10061) );
  nd02d1 U7568 ( .A1(n8831), .A2(n6892), .ZN(n10282) );
  inv0d0 U7569 ( .I(n8935), .ZN(n2792) );
  inv0d0 U7570 ( .I(n8675), .ZN(n3036) );
  nd02d1 U7571 ( .A1(N13666), .A2(n11997), .ZN(n8621) );
  nr02d1 U7572 ( .A1(n8091), .A2(n7081), .ZN(n5777) );
  inv0d0 U7575 ( .I(n7530), .ZN(n4185) );
  nr02d1 U7576 ( .A1(n11457), .A2(n7097), .ZN(n11454) );
  nr13d1 U7577 ( .A1(N8549), .A2(n8208), .A3(n8957), .ZN(n8956) );
  inv0d0 U7578 ( .I(n5251), .ZN(n3896) );
  nr02d1 U7579 ( .A1(n5261), .A2(n5262), .ZN(n5260) );
  inv0d0 U7580 ( .I(n2424), .ZN(n2427) );
  inv0d0 U7581 ( .I(n10378), .ZN(n3092) );
  inv0d0 U7582 ( .I(n8574), .ZN(n3352) );
  inv0d0 U7583 ( .I(n8579), .ZN(n3390) );
  inv0d0 U7584 ( .I(n5117), .ZN(n3908) );
  nd03d1 U7585 ( .A1(n5201), .A2(n4698), .A3(N10701), .ZN(n6030) );
  nr02d1 U7587 ( .A1(n4791), .A2(n9504), .ZN(n8041) );
  inv0d0 U7588 ( .I(n6208), .ZN(n3356) );
  aoim22d1 U7590 ( .A1(n6111), .A2(n7010), .B1(n7011), .B2(n7012), .Z(n7009)
         );
  nr02d1 U7591 ( .A1(n4675), .A2(n5388), .ZN(n6167) );
  nr02d1 U7592 ( .A1(n9975), .A2(n7410), .ZN(n9974) );
  inv0d0 U7593 ( .I(n9980), .ZN(n3505) );
  nr02d1 U7597 ( .A1(n7442), .A2(n8290), .ZN(n12064) );
  nr02d1 U7599 ( .A1(n11323), .A2(n9671), .ZN(n7472) );
  inv0d0 U7600 ( .I(n8055), .ZN(n3049) );
  nd02d1 U7601 ( .A1(n12040), .A2(n5745), .ZN(n4456) );
  nr02d1 U7602 ( .A1(n6817), .A2(n10297), .ZN(n11932) );
  nd02d1 U7604 ( .A1(N12098), .A2(n4484), .ZN(n5382) );
  nr02d1 U7605 ( .A1(n11878), .A2(n10368), .ZN(n11970) );
  nr02d1 U7609 ( .A1(n8801), .A2(n7340), .ZN(n8800) );
  aoi31d1 U7610 ( .B1(n1294), .B2(n1237), .B3(n2068), .A(n1330), .ZN(n26) );
  nr02d1 U7611 ( .A1(n5235), .A2(n11980), .ZN(n10172) );
  nr02d1 U7614 ( .A1(n7396), .A2(n7400), .ZN(n5731) );
  nr02d1 U7615 ( .A1(n7375), .A2(n6415), .ZN(n4961) );
  nr02d1 U7616 ( .A1(n4277), .A2(n6685), .ZN(n11342) );
  inv0d0 U7619 ( .I(n8084), .ZN(n3847) );
  nr02d1 U7621 ( .A1(n5834), .A2(n12030), .ZN(n12032) );
  inv0d0 U7622 ( .I(n7605), .ZN(n4129) );
  nr02d1 U7625 ( .A1(n6166), .A2(n3268), .ZN(n6277) );
  nr02d1 U7627 ( .A1(n6088), .A2(n10726), .ZN(n8440) );
  nr02d1 U7630 ( .A1(n6051), .A2(n6397), .ZN(n8870) );
  nr02d1 U7631 ( .A1(n4483), .A2(n5265), .ZN(n4485) );
  nr02d1 U7635 ( .A1(n6998), .A2(n5825), .ZN(n5721) );
  nr02d1 U7636 ( .A1(n7205), .A2(n6084), .ZN(n4956) );
  nd02d1 U7640 ( .A1(n11673), .A2(n3438), .ZN(n6181) );
  nd02d1 U7641 ( .A1(N12498), .A2(n11680), .ZN(n9315) );
  nr02d1 U7642 ( .A1(n8888), .A2(n11325), .ZN(n11324) );
  nr02d1 U7643 ( .A1(n6597), .A2(n10931), .ZN(n8069) );
  nd02d1 U7646 ( .A1(N12066), .A2(n7046), .ZN(n9273) );
  nd02d1 U7647 ( .A1(N12658), .A2(n11696), .ZN(n4538) );
  nd02d1 U7648 ( .A1(N13394), .A2(n5488), .ZN(n5491) );
  nr02d1 U7649 ( .A1(n6619), .A2(n5308), .ZN(n5751) );
  inv0d0 U7650 ( .I(n10791), .ZN(n3582) );
  nr02d1 U7651 ( .A1(n8445), .A2(n10726), .ZN(n5309) );
  inv0d0 U7656 ( .I(n5576), .ZN(n3026) );
  nr02d1 U7657 ( .A1(n11180), .A2(n8020), .ZN(n11951) );
  nd02d1 U7659 ( .A1(n5201), .A2(n5765), .ZN(n6028) );
  nr02d1 U7660 ( .A1(n10357), .A2(n8781), .ZN(n7356) );
  inv0d0 U7662 ( .I(n8670), .ZN(n3225) );
  nd02d1 U7663 ( .A1(N9106), .A2(n5456), .ZN(n11425) );
  inv0d0 U7664 ( .I(n8113), .ZN(n4289) );
  nd02d1 U7665 ( .A1(n8401), .A2(n7685), .ZN(n5216) );
  inv0d0 U7668 ( .I(n8765), .ZN(n2996) );
  inv0d0 U7670 ( .I(n9617), .ZN(n3547) );
  inv0d0 U7672 ( .I(n6181), .ZN(n3437) );
  inv0d0 U7675 ( .I(n8497), .ZN(n3552) );
  nr02d1 U7676 ( .A1(n6855), .A2(n10722), .ZN(n11605) );
  nr02d1 U7677 ( .A1(n11242), .A2(n9312), .ZN(n10844) );
  nr02d1 U7680 ( .A1(n5798), .A2(n7332), .ZN(n11968) );
  nr02d1 U7682 ( .A1(n5053), .A2(n6843), .ZN(n6845) );
  nr02d1 U7683 ( .A1(n3800), .A2(n7076), .ZN(n9952) );
  nd03d1 U7684 ( .A1(n7444), .A2(n5458), .A3(n8264), .ZN(n8272) );
  nr02d1 U7688 ( .A1(n6123), .A2(n7645), .ZN(n8869) );
  nr02d1 U7692 ( .A1(n8796), .A2(n10279), .ZN(n6549) );
  inv0d0 U7693 ( .I(n7298), .ZN(n2921) );
  nr02d1 U7697 ( .A1(n3302), .A2(n6997), .ZN(n10951) );
  inv0d0 U7698 ( .I(n4631), .ZN(n3296) );
  nr02d1 U7705 ( .A1(n4955), .A2(n4712), .ZN(n4714) );
  nr02d1 U7706 ( .A1(n6337), .A2(n4969), .ZN(n6351) );
  inv0d0 U7707 ( .I(n9406), .ZN(n3263) );
  nr02d1 U7709 ( .A1(n8579), .A2(n8570), .ZN(n5464) );
  nr02d1 U7710 ( .A1(n5853), .A2(n6768), .ZN(n5025) );
  nr02d1 U7711 ( .A1(n6368), .A2(n9379), .ZN(n4592) );
  nr02d1 U7713 ( .A1(n5859), .A2(n9769), .ZN(n8266) );
  nr02d1 U7714 ( .A1(n6805), .A2(n6764), .ZN(n9018) );
  nr02d1 U7715 ( .A1(n6740), .A2(n8222), .ZN(n7453) );
  nr02d1 U7716 ( .A1(n6759), .A2(n5321), .ZN(n11615) );
  nr02d1 U7719 ( .A1(n6655), .A2(n5322), .ZN(n8782) );
  nd02d1 U7720 ( .A1(n3281), .A2(n4419), .ZN(n6311) );
  nr02d1 U7721 ( .A1(n4139), .A2(n8107), .ZN(n7444) );
  nr02d1 U7722 ( .A1(n5359), .A2(n5358), .ZN(n8486) );
  nd02d1 U7726 ( .A1(n9276), .A2(n3425), .ZN(n4478) );
  nr02d1 U7730 ( .A1(n4765), .A2(n4942), .ZN(n4784) );
  nd02d1 U7731 ( .A1(N13554), .A2(n6340), .ZN(n6353) );
  nr02d1 U7732 ( .A1(n11933), .A2(n4919), .ZN(n11935) );
  nr02d1 U7733 ( .A1(n6529), .A2(n5046), .ZN(n6243) );
  nd02d1 U7734 ( .A1(n8508), .A2(n5642), .ZN(n8520) );
  nd02d1 U7739 ( .A1(n8039), .A2(n8045), .ZN(n5698) );
  nd03d1 U7740 ( .A1(n6232), .A2(n5927), .A3(n3402), .ZN(n12013) );
  nd03d1 U7741 ( .A1(n5140), .A2(n4950), .A3(n6451), .ZN(n6470) );
  aoim22d1 U7742 ( .A1(n2826), .A2(n11118), .B1(n11119), .B2(n4929), .Z(n11115) );
  nr02d1 U7744 ( .A1(n5030), .A2(n6830), .ZN(n9073) );
  nr02d1 U7745 ( .A1(n3465), .A2(n7150), .ZN(n10019) );
  inv0d0 U7746 ( .I(n7690), .ZN(n3877) );
  nr02d1 U7747 ( .A1(n5218), .A2(n9163), .ZN(n9170) );
  nr02d1 U7748 ( .A1(n5535), .A2(n6183), .ZN(n11681) );
  nd02d1 U7751 ( .A1(N14322), .A2(n6456), .ZN(n8695) );
  nd02d1 U7753 ( .A1(n8433), .A2(n6931), .ZN(n10707) );
  nd02d1 U7754 ( .A1(N13074), .A2(n6271), .ZN(n6281) );
  nd02d1 U7755 ( .A1(n3785), .A2(n5337), .ZN(n7011) );
  nd02d1 U7759 ( .A1(N13746), .A2(n11991), .ZN(n10126) );
  inv0d0 U7760 ( .I(n6334), .ZN(n2802) );
  inv0d0 U7761 ( .I(n6000), .ZN(n3975) );
  nr02d1 U7762 ( .A1(n6259), .A2(n6631), .ZN(n6629) );
  nr02d1 U7764 ( .A1(n5379), .A2(n4478), .ZN(n5378) );
  nd02d1 U7766 ( .A1(N13250), .A2(n12000), .ZN(n7385) );
  inv0d0 U7767 ( .I(n7431), .ZN(n3901) );
  nr02d1 U7768 ( .A1(n7266), .A2(n4955), .ZN(n7270) );
  inv0d0 U7771 ( .I(n7610), .ZN(n3989) );
  inv0d0 U7772 ( .I(n4585), .ZN(n3322) );
  nr02d1 U7773 ( .A1(n6988), .A2(n6987), .ZN(n7724) );
  nr02d1 U7778 ( .A1(n6658), .A2(n6492), .ZN(n8730) );
  nr02d1 U7779 ( .A1(n6059), .A2(n5270), .ZN(n9189) );
  nd03d1 U7782 ( .A1(n3530), .A2(n8471), .A3(n3534), .ZN(n6128) );
  nr02d1 U7784 ( .A1(n9757), .A2(n5958), .ZN(n9758) );
  nr02d1 U7786 ( .A1(n8829), .A2(n11960), .ZN(n4925) );
  inv0d0 U7789 ( .I(n8798), .ZN(n2865) );
  nd02d1 U7791 ( .A1(N8471), .A2(n10426), .ZN(n6711) );
  inv0d0 U7794 ( .I(n2601), .ZN(N8471) );
  inv0d0 U7796 ( .I(n2600), .ZN(n2602) );
  nr02d1 U7797 ( .A1(n6529), .A2(n5397), .ZN(n5722) );
  nr02d1 U7798 ( .A1(n2999), .A2(n4817), .ZN(n5651) );
  nr02d1 U7801 ( .A1(n6736), .A2(n10988), .ZN(n10991) );
  nr02d1 U7802 ( .A1(n4953), .A2(n4722), .ZN(n4723) );
  inv0d0 U7803 ( .I(n8179), .ZN(n4278) );
  nd02d1 U7804 ( .A1(n9076), .A2(n5855), .ZN(n7439) );
  nd02d1 U7806 ( .A1(n4804), .A2(n2955), .ZN(n4807) );
  nr02d1 U7807 ( .A1(n9066), .A2(n8873), .ZN(n6815) );
  nr02d1 U7808 ( .A1(n10661), .A2(n6927), .ZN(n9144) );
  inv0d0 U7813 ( .I(n6485), .ZN(n3107) );
  inv0d0 U7816 ( .I(n6477), .ZN(n3131) );
  nr02d1 U7817 ( .A1(n10952), .A2(n3306), .ZN(n5719) );
  inv0d0 U7818 ( .I(n10953), .ZN(n3306) );
  nr02d1 U7819 ( .A1(n6402), .A2(n4963), .ZN(n5711) );
  aoim22d1 U7821 ( .A1(n3295), .A2(n10949), .B1(n9404), .B2(n10950), .Z(n10938) );
  inv0d0 U7822 ( .I(n9401), .ZN(n3295) );
  nr02d1 U7823 ( .A1(n7504), .A2(n7457), .ZN(n7505) );
  inv0d0 U7824 ( .I(n11427), .ZN(n4144) );
  nr02d1 U7826 ( .A1(n8968), .A2(n5862), .ZN(n8973) );
  nd02d1 U7828 ( .A1(N9596), .A2(n11470), .ZN(n6835) );
  inv0d0 U7829 ( .I(n5170), .ZN(n3940) );
  nd02d1 U7830 ( .A1(N12818), .A2(n12012), .ZN(n9346) );
  nd02d1 U7832 ( .A1(n4047), .A2(n11271), .ZN(n4389) );
  nr02d1 U7836 ( .A1(n8416), .A2(n5262), .ZN(n4412) );
  nr02d1 U7837 ( .A1(n7469), .A2(n4342), .ZN(n7477) );
  nd03d1 U7839 ( .A1(n8045), .A2(n3008), .A3(N14722), .ZN(n9504) );
  inv0d0 U7843 ( .I(n6281), .ZN(n3270) );
  aoim22d1 U7850 ( .A1(n4046), .A2(n9838), .B1(n9839), .B2(n9840), .Z(n9837)
         );
  inv0d0 U7851 ( .I(n6407), .ZN(n3236) );
  nr02d1 U7852 ( .A1(n8334), .A2(n7640), .ZN(n8336) );
  inv0d0 U7853 ( .I(n9853), .ZN(n3902) );
  aoim22d1 U7857 ( .A1(n9255), .A2(n10396), .B1(n9261), .B2(n10395), .Z(n9993)
         );
  inv0d0 U7858 ( .I(n9616), .ZN(n3490) );
  nd02d1 U7860 ( .A1(N12786), .A2(n12009), .ZN(n7132) );
  inv0d0 U7865 ( .I(n7735), .ZN(n3776) );
  nr02d1 U7866 ( .A1(n7166), .A2(n7433), .ZN(n8866) );
  nr02d1 U7868 ( .A1(n3328), .A2(n5732), .ZN(n12001) );
  nr02d1 U7872 ( .A1(n6346), .A2(n3303), .ZN(n5718) );
  inv0d0 U7875 ( .I(n6333), .ZN(n3303) );
  nd02d1 U7876 ( .A1(N13794), .A2(n11989), .ZN(n6380) );
  nr02d1 U7877 ( .A1(n8074), .A2(n8546), .ZN(n8542) );
  nd02d1 U7881 ( .A1(N12802), .A2(n9610), .ZN(n9342) );
  inv0d0 U7882 ( .I(n6648), .ZN(n4009) );
  inv0d0 U7883 ( .I(n7000), .ZN(n2803) );
  inv0d0 U7885 ( .I(n7241), .ZN(n3198) );
  nr02d1 U7886 ( .A1(n6504), .A2(n5698), .ZN(n6514) );
  inv0d0 U7888 ( .I(n8449), .ZN(n3766) );
  inv0d0 U7891 ( .I(n7740), .ZN(n3786) );
  nr02d1 U7892 ( .A1(n4963), .A2(n4670), .ZN(n4674) );
  nd02d1 U7893 ( .A1(n8268), .A2(n6496), .ZN(n5876) );
  inv0d0 U7895 ( .I(n5884), .ZN(n4062) );
  aoim22d1 U7897 ( .A1(n2943), .A2(n6513), .B1(n6514), .B2(n5639), .Z(n6511)
         );
  inv0d0 U7898 ( .I(n5641), .ZN(n2943) );
  nd02d1 U7899 ( .A1(n7128), .A2(n10883), .ZN(n8850) );
  aoim22d1 U7901 ( .A1(n7715), .A2(n6073), .B1(n7714), .B2(n5268), .Z(n7713)
         );
  nd02d1 U7902 ( .A1(n10480), .A2(n10489), .ZN(n7458) );
  nd02d1 U7904 ( .A1(n7761), .A2(n5001), .ZN(n7769) );
  nr02d1 U7905 ( .A1(n11496), .A2(n5786), .ZN(n11498) );
  inv0d0 U7908 ( .I(n5708), .ZN(n4901) );
  inv0d0 U7910 ( .I(n9073), .ZN(n4089) );
  nr02d1 U7911 ( .A1(n7087), .A2(n7072), .ZN(n11677) );
  inv0d0 U7914 ( .I(n6306), .ZN(n3315) );
  nd03d1 U7915 ( .A1(n4102), .A2(n6547), .A3(N9498), .ZN(n9071) );
  nd02d1 U7916 ( .A1(n11191), .A2(n2862), .ZN(n8801) );
  nd02d1 U7917 ( .A1(N14130), .A2(n11981), .ZN(n7919) );
  nr13d1 U7918 ( .A1(N9260), .A2(n10555), .A3(n5284), .ZN(n5886) );
  nr02d1 U7919 ( .A1(n5920), .A2(n6318), .ZN(n8070) );
  nd02d1 U7920 ( .A1(n6688), .A2(n8119), .ZN(n6694) );
  nr02d1 U7921 ( .A1(n4255), .A2(n8214), .ZN(n7454) );
  nr02d1 U7922 ( .A1(n6893), .A2(n5135), .ZN(n8867) );
  nr02d1 U7923 ( .A1(n6562), .A2(n5156), .ZN(n5725) );
  inv0d0 U7925 ( .I(n8410), .ZN(n3875) );
  nr02d1 U7929 ( .A1(n8574), .A2(n4982), .ZN(n8580) );
  nr02d1 U7930 ( .A1(n5268), .A2(n10707), .ZN(n6976) );
  nr02d1 U7931 ( .A1(n4959), .A2(n6693), .ZN(n9846) );
  nd02d1 U7932 ( .A1(n8852), .A2(n3410), .ZN(n6216) );
  nr02d1 U7937 ( .A1(n7604), .A2(n6363), .ZN(n7217) );
  nd03d1 U7939 ( .A1(n3533), .A2(n8471), .A3(n3532), .ZN(n9981) );
  nr02d1 U7940 ( .A1(n6565), .A2(n5164), .ZN(n8524) );
  nd02d1 U7942 ( .A1(n8238), .A2(n6666), .ZN(n8243) );
  nr02d1 U7944 ( .A1(n4663), .A2(n10861), .ZN(n12016) );
  nd02d1 U7945 ( .A1(n3012), .A2(n8738), .ZN(n9500) );
  nd02d1 U7946 ( .A1(n6026), .A2(n5765), .ZN(n6035) );
  nr02d1 U7947 ( .A1(n6065), .A2(n5755), .ZN(n6068) );
  nd02d1 U7948 ( .A1(n10400), .A2(n3539), .ZN(n7760) );
  nr02d1 U7949 ( .A1(n6397), .A2(n11484), .ZN(n8317) );
  nr02d1 U7950 ( .A1(n11448), .A2(n5918), .ZN(n11450) );
  nd02d1 U7951 ( .A1(n11710), .A2(n3372), .ZN(n10393) );
  nr02d1 U7952 ( .A1(n11689), .A2(n6188), .ZN(n4522) );
  nr02d1 U7953 ( .A1(n7222), .A2(n7147), .ZN(n12002) );
  nr02d1 U7954 ( .A1(n5988), .A2(n3317), .ZN(n10918) );
  nr02d1 U7956 ( .A1(n4918), .A2(n4919), .ZN(n4897) );
  nd02d1 U7957 ( .A1(N12994), .A2(n12005), .ZN(n5462) );
  nr02d1 U7958 ( .A1(n6366), .A2(n9422), .ZN(n8624) );
  nr02d1 U7961 ( .A1(n6391), .A2(n10984), .ZN(n7230) );
  nr02d1 U7962 ( .A1(n7848), .A2(n6294), .ZN(n7853) );
  nr02d1 U7963 ( .A1(n6641), .A2(n5809), .ZN(n11392) );
  nr02d1 U7964 ( .A1(n5600), .A2(n11047), .ZN(n7956) );
  nd02d1 U7965 ( .A1(n11992), .A2(n9425), .ZN(n8626) );
  nd12d1 U7966 ( .A1(n1861), .A2(n11709), .ZN(n7125) );
  nd12d1 U7967 ( .A1(n9461), .A2(n9459), .ZN(n4729) );
  inv0d0 U7969 ( .I(n7410), .ZN(n3524) );
  nr02d1 U7970 ( .A1(n10164), .A2(n5235), .ZN(n10173) );
  nd02d1 U7971 ( .A1(N12050), .A2(n5377), .ZN(n5379) );
  nr02d1 U7972 ( .A1(n5074), .A2(n4491), .ZN(n5070) );
  nr02d1 U7973 ( .A1(n4947), .A2(n4999), .ZN(n5701) );
  nd02d1 U7974 ( .A1(n4946), .A2(n6466), .ZN(n6158) );
  nr02d1 U7975 ( .A1(n4483), .A2(n7237), .ZN(n8075) );
  nd02d1 U7978 ( .A1(n8434), .A2(n5655), .ZN(n8437) );
  inv0d0 U7979 ( .I(n2523), .ZN(N8868) );
  inv0d0 U7983 ( .I(n8072), .ZN(n3266) );
  nd03d1 U7984 ( .A1(n3807), .A2(n7153), .A3(N11226), .ZN(n6985) );
  inv0d0 U7985 ( .I(n2086), .ZN(n2088) );
  nr02d1 U7987 ( .A1(n7955), .A2(n11047), .ZN(n11840) );
  nd03d1 U7990 ( .A1(n11087), .A2(n5979), .A3(n8047), .ZN(n9511) );
  nr02d1 U7991 ( .A1(n6919), .A2(n5737), .ZN(n6603) );
  nr02d1 U7992 ( .A1(n6151), .A2(n11244), .ZN(n5367) );
  nr02d1 U7993 ( .A1(n11838), .A2(n6564), .ZN(n11839) );
  inv0d0 U7994 ( .I(n9612), .ZN(n3340) );
  nd02d1 U7997 ( .A1(N12754), .A2(n8852), .ZN(n6226) );
  nr02d1 U7999 ( .A1(n9312), .A2(n3442), .ZN(n10039) );
  nd03d1 U8000 ( .A1(n7455), .A2(n4331), .A3(n4269), .ZN(n11373) );
  nr02d1 U8001 ( .A1(n6987), .A2(n6088), .ZN(n9626) );
  nd02d1 U8002 ( .A1(n5213), .A2(n10426), .ZN(n12072) );
  nd03d1 U8003 ( .A1(n7456), .A2(n6719), .A3(n11356), .ZN(n11367) );
  nr02d1 U8004 ( .A1(n6643), .A2(n10609), .ZN(n5081) );
  nr02d1 U8007 ( .A1(n5246), .A2(n3856), .ZN(n6046) );
  nr02d1 U8009 ( .A1(n4300), .A2(n11053), .ZN(n11978) );
  nd03d1 U8010 ( .A1(n11673), .A2(n3438), .A3(n3436), .ZN(n5403) );
  nr02d1 U8012 ( .A1(n7349), .A2(n7350), .ZN(n4864) );
  nd03d1 U8013 ( .A1(n6652), .A2(n5579), .A3(n7584), .ZN(n7592) );
  nr02d1 U8014 ( .A1(n5684), .A2(n7619), .ZN(n12063) );
  nd02d1 U8015 ( .A1(n8654), .A2(n5364), .ZN(n8664) );
  nd02d1 U8016 ( .A1(N9064), .A2(n11286), .ZN(n5016) );
  nd02d1 U8019 ( .A1(n8984), .A2(n4205), .ZN(n8989) );
  nr02d1 U8022 ( .A1(n6356), .A2(n4633), .ZN(n7341) );
  nr02d1 U8023 ( .A1(n8909), .A2(n10459), .ZN(n7468) );
  nr02d1 U8024 ( .A1(n5774), .A2(n5846), .ZN(n8865) );
  nr02d1 U8028 ( .A1(n7123), .A2(n8563), .ZN(n8848) );
  nd02d1 U8029 ( .A1(n11919), .A2(n4924), .ZN(n4885) );
  nr02d1 U8033 ( .A1(n4756), .A2(n7955), .ZN(n8718) );
  nr02d1 U8034 ( .A1(n10389), .A2(n6394), .ZN(n11983) );
  inv0d0 U8035 ( .I(n7836), .ZN(n2798) );
  nr02d1 U8036 ( .A1(n9679), .A2(n11330), .ZN(n11297) );
  nr02d1 U8037 ( .A1(n4419), .A2(n6313), .ZN(n11753) );
  nr02d1 U8040 ( .A1(n5698), .A2(n4942), .ZN(n11861) );
  nr02d1 U8042 ( .A1(n5709), .A2(n6993), .ZN(n6579) );
  nr02d1 U8045 ( .A1(n6927), .A2(n8380), .ZN(n6926) );
  inv0d0 U8047 ( .I(n6062), .ZN(n3723) );
  inv0d0 U8049 ( .I(n7561), .ZN(n4169) );
  aoim22d1 U8050 ( .A1(n11682), .A2(n3447), .B1(n4515), .B2(n3495), .Z(n11674)
         );
  inv0d0 U8051 ( .I(n11685), .ZN(n3495) );
  nr02d1 U8052 ( .A1(n3500), .A2(n4515), .ZN(n4513) );
  inv0d0 U8053 ( .I(n6076), .ZN(n3753) );
  inv0d0 U8054 ( .I(n6725), .ZN(n4263) );
  nr02d1 U8056 ( .A1(n6091), .A2(n6619), .ZN(n6102) );
  inv0d0 U8057 ( .I(n8414), .ZN(n3895) );
  nr02d1 U8058 ( .A1(n9691), .A2(n8126), .ZN(n8930) );
  nd03d1 U8060 ( .A1(n7456), .A2(n6719), .A3(n6709), .ZN(n6722) );
  inv0d0 U8063 ( .I(n5616), .ZN(n3088) );
  nr02d1 U8065 ( .A1(n6358), .A2(n4635), .ZN(n9510) );
  inv0d0 U8067 ( .I(n4714), .ZN(n3021) );
  nr02d1 U8068 ( .A1(n9590), .A2(n11130), .ZN(n11965) );
  nr02d1 U8069 ( .A1(n8357), .A2(n8091), .ZN(n8364) );
  inv0d0 U8070 ( .I(n11407), .ZN(n4510) );
  nr02d1 U8071 ( .A1(n6066), .A2(n5280), .ZN(n6969) );
  nr02d1 U8073 ( .A1(n10983), .A2(n6291), .ZN(n11221) );
  nr02d1 U8074 ( .A1(n5879), .A2(n6138), .ZN(n9037) );
  nr02d1 U8078 ( .A1(n10047), .A2(n6098), .ZN(n10051) );
  nr02d1 U8079 ( .A1(n10735), .A2(n11613), .ZN(n7736) );
  nr02d1 U8080 ( .A1(n9361), .A2(n5825), .ZN(n9372) );
  inv0d0 U8081 ( .I(n7458), .ZN(n4244) );
  nd03d1 U8082 ( .A1(N9092), .A2(n11423), .A3(n4172), .ZN(n5861) );
  nr02d1 U8085 ( .A1(n6150), .A2(n6612), .ZN(n6609) );
  inv0d0 U8086 ( .I(n5040), .ZN(n4096) );
  nr13d1 U8087 ( .A1(N9951), .A2(n9836), .A3(n5098), .ZN(n5088) );
  nr13d1 U8088 ( .A1(n7035), .A2(n7036), .A3(n7037), .ZN(n7032) );
  inv0d0 U8091 ( .I(n8077), .ZN(n3572) );
  nd03d1 U8092 ( .A1(n9726), .A2(n11372), .A3(n8967), .ZN(n8215) );
  nr13d1 U8093 ( .A1(n5752), .A2(n5294), .A3(n5296), .ZN(n5304) );
  nd03d1 U8094 ( .A1(n9072), .A2(n4102), .A3(N9512), .ZN(n5940) );
  nd02d1 U8095 ( .A1(n7515), .A2(n8118), .ZN(n7512) );
  inv0d0 U8097 ( .I(n11508), .ZN(n3992) );
  nr02d1 U8101 ( .A1(n4689), .A2(n6618), .ZN(n9621) );
  nr02d1 U8102 ( .A1(n6330), .A2(n11274), .ZN(n10608) );
  inv0d0 U8103 ( .I(n6667), .ZN(n4157) );
  inv0d0 U8104 ( .I(n1221), .ZN(n1269) );
  nr02d1 U8105 ( .A1(n8172), .A2(n6146), .ZN(n8177) );
  inv0d0 U8106 ( .I(n4952), .ZN(n3053) );
  inv0d0 U8107 ( .I(n9062), .ZN(n4076) );
  nr02d1 U8114 ( .A1(n7812), .A2(n7811), .ZN(n4525) );
  nr02d1 U8115 ( .A1(n10762), .A2(n8464), .ZN(n11637) );
  inv0d0 U8116 ( .I(n5350), .ZN(n4949) );
  nr02d1 U8117 ( .A1(n9625), .A2(n9201), .ZN(n9212) );
  nr02d1 U8119 ( .A1(n8222), .A2(n4222), .ZN(n8225) );
  nd03d1 U8120 ( .A1(n8894), .A2(n4858), .A3(N8044), .ZN(n8130) );
  inv0d0 U8121 ( .I(n8679), .ZN(n3128) );
  inv0d0 U8122 ( .I(n5823), .ZN(n4150) );
  nd02d1 U8126 ( .A1(N8562), .A2(n6720), .ZN(n11362) );
  nr02d1 U8127 ( .A1(n5607), .A2(n7117), .ZN(n8751) );
  nd03d1 U8128 ( .A1(n3471), .A2(n6167), .A3(n6168), .ZN(n6164) );
  inv0d0 U8129 ( .I(n7724), .ZN(n3803) );
  nd02d1 U8130 ( .A1(n8127), .A2(n11333), .ZN(n9688) );
  nd02d1 U8131 ( .A1(n8967), .A2(n11372), .ZN(n8974) );
  nr02d1 U8132 ( .A1(n4963), .A2(n6399), .ZN(n6398) );
  nd02d1 U8133 ( .A1(n7128), .A2(n7137), .ZN(n10883) );
  nr02d1 U8134 ( .A1(n6735), .A2(n7452), .ZN(n6743) );
  inv0d0 U8136 ( .I(n5716), .ZN(n5044) );
  nd03d1 U8137 ( .A1(n4176), .A2(n11286), .A3(n5025), .ZN(n8259) );
  inv0d0 U8141 ( .I(n5499), .ZN(n2808) );
  nd02d1 U8145 ( .A1(n10203), .A2(n5354), .ZN(n6492) );
  nd02d1 U8148 ( .A1(n5170), .A2(n6003), .ZN(n6002) );
  nr02d1 U8149 ( .A1(n8107), .A2(n7447), .ZN(n6660) );
  nr02d1 U8151 ( .A1(n11828), .A2(n7948), .ZN(n11830) );
  nr02d1 U8155 ( .A1(n4395), .A2(n11253), .ZN(n7751) );
  inv0d0 U8156 ( .I(n7954), .ZN(n5140) );
  nr02d1 U8157 ( .A1(n5927), .A2(n8563), .ZN(n12010) );
  nd02d1 U8158 ( .A1(n5780), .A2(n6870), .ZN(n6876) );
  inv0d0 U8161 ( .I(n6650), .ZN(n4966) );
  nr02d1 U8162 ( .A1(n11802), .A2(n7375), .ZN(n11808) );
  inv0d0 U8163 ( .I(n6595), .ZN(n5380) );
  nd03d1 U8168 ( .A1(n6478), .A2(n4300), .A3(n9599), .ZN(n8052) );
  nd02d1 U8169 ( .A1(n9429), .A2(n4416), .ZN(n7882) );
  inv0d0 U8170 ( .I(n9501), .ZN(n3008) );
  nd03d1 U8171 ( .A1(n4559), .A2(n6253), .A3(n9355), .ZN(n9354) );
  inv0d0 U8174 ( .I(n7822), .ZN(n2797) );
  nd02d1 U8177 ( .A1(n6456), .A2(n6556), .ZN(n10384) );
  inv0d0 U8178 ( .I(n8744), .ZN(n2937) );
  nd03d1 U8180 ( .A1(n11083), .A2(n8043), .A3(n8041), .ZN(n11082) );
  nd02d1 U8181 ( .A1(N12978), .A2(n11723), .ZN(n11721) );
  nr02d1 U8182 ( .A1(n7357), .A2(n9525), .ZN(n8772) );
  inv0d0 U8183 ( .I(n6573), .ZN(n4411) );
  nr02d1 U8184 ( .A1(n5766), .A2(n5196), .ZN(n5199) );
  inv0d0 U8185 ( .I(n5807), .ZN(n5778) );
  nr02d1 U8186 ( .A1(n5596), .A2(n5702), .ZN(n5603) );
  inv0d0 U8188 ( .I(n6960), .ZN(n3870) );
  inv0d0 U8193 ( .I(n10746), .ZN(n3780) );
  nr13d1 U8194 ( .A1(n6111), .A2(n10745), .A3(n10746), .ZN(n10744) );
  nr02d1 U8195 ( .A1(n10366), .A2(n10368), .ZN(n11971) );
  nd03d1 U8197 ( .A1(n8695), .A2(n5136), .A3(n3123), .ZN(n7364) );
  nd02d1 U8200 ( .A1(n12001), .A2(n6908), .ZN(n9376) );
  nd02d1 U8201 ( .A1(N11778), .A2(n12040), .ZN(n9989) );
  inv0d0 U8202 ( .I(n6409), .ZN(n3239) );
  nd02d1 U8203 ( .A1(n8118), .A2(n6720), .ZN(n10500) );
  inv0d0 U8204 ( .I(n8644), .ZN(n3235) );
  nr02d1 U8205 ( .A1(n8664), .A2(n5708), .ZN(n8668) );
  nr02d1 U8206 ( .A1(n10396), .A2(n5834), .ZN(n10395) );
  nr02d1 U8208 ( .A1(n5396), .A2(n10823), .ZN(n4498) );
  inv0d0 U8209 ( .I(n5392), .ZN(n3471) );
  nd02d1 U8213 ( .A1(n7814), .A2(n7391), .ZN(n7816) );
  inv0d0 U8214 ( .I(n7411), .ZN(n5427) );
  nr02d1 U8216 ( .A1(n5807), .A2(n6743), .ZN(n6746) );
  inv0d0 U8222 ( .I(n5262), .ZN(n3858) );
  nr02d1 U8224 ( .A1(n9331), .A2(n4990), .ZN(n9337) );
  nd03d1 U8226 ( .A1(n7952), .A2(n5136), .A3(n3123), .ZN(n11033) );
  inv0d0 U8228 ( .I(n9012), .ZN(n4152) );
  inv0d0 U8229 ( .I(n5709), .ZN(n5364) );
  nr02d1 U8230 ( .A1(n6098), .A2(n11689), .ZN(n12018) );
  nr02d1 U8231 ( .A1(n6885), .A2(n6039), .ZN(n6888) );
  nr02d1 U8232 ( .A1(n3214), .A2(n4694), .ZN(n5557) );
  nr02d1 U8233 ( .A1(n9536), .A2(n11196), .ZN(n8785) );
  nr02d1 U8234 ( .A1(n6242), .A2(n4311), .ZN(n9619) );
  nr02d1 U8235 ( .A1(n5737), .A2(n7232), .ZN(n9613) );
  nr02d1 U8237 ( .A1(n5600), .A2(n11840), .ZN(n7957) );
  nd02d1 U8238 ( .A1(n9023), .A2(n4323), .ZN(n9027) );
  inv0d0 U8239 ( .I(n11130), .ZN(n2864) );
  nr02d1 U8240 ( .A1(n6371), .A2(n10058), .ZN(n10060) );
  inv0d0 U8241 ( .I(n11849), .ZN(n3010) );
  nr02d1 U8242 ( .A1(n6970), .A2(n5755), .ZN(n6973) );
  nd02d1 U8244 ( .A1(n4914), .A2(n11953), .ZN(n11180) );
  nr02d1 U8245 ( .A1(n8520), .A2(n5733), .ZN(n8525) );
  nd02d1 U8247 ( .A1(n8936), .A2(n6697), .ZN(n8945) );
  nd02d1 U8248 ( .A1(n8567), .A2(n7388), .ZN(n8574) );
  nr02d1 U8249 ( .A1(n11627), .A2(n6113), .ZN(n11629) );
  nd03d1 U8250 ( .A1(n10386), .A2(n5728), .A3(n3043), .ZN(n4708) );
  nd02d1 U8251 ( .A1(n10676), .A2(n3832), .ZN(n5198) );
  inv0d0 U8255 ( .I(n6983), .ZN(n3650) );
  nr02d1 U8258 ( .A1(n11588), .A2(n6622), .ZN(n11589) );
  nd02d1 U8259 ( .A1(n9032), .A2(n4118), .ZN(n5874) );
  nr02d1 U8260 ( .A1(n6371), .A2(n3412), .ZN(n12017) );
  nd02d1 U8261 ( .A1(n8452), .A2(n5427), .ZN(n8455) );
  nr02d1 U8263 ( .A1(n5249), .A2(n9376), .ZN(n11741) );
  inv0d0 U8264 ( .I(n7657), .ZN(n3976) );
  nd02d1 U8265 ( .A1(N13442), .A2(n8601), .ZN(n11770) );
  nd02d1 U8268 ( .A1(n3330), .A2(n5732), .ZN(n6283) );
  inv0d0 U8269 ( .I(n5926), .ZN(n5579) );
  nd02d1 U8271 ( .A1(N13826), .A2(n9429), .ZN(n7884) );
  inv0d0 U8273 ( .I(n5994), .ZN(n3963) );
  nd02d1 U8276 ( .A1(n5259), .A2(n4477), .ZN(n4490) );
  nd02d1 U8277 ( .A1(N8666), .A2(n12071), .ZN(n8971) );
  nd02d1 U8278 ( .A1(n10969), .A2(n6600), .ZN(n7223) );
  inv0d0 U8279 ( .I(n6812), .ZN(n4102) );
  nd02d1 U8280 ( .A1(n10795), .A2(n4946), .ZN(n12026) );
  nd02d1 U8282 ( .A1(n10468), .A2(n4292), .ZN(n8176) );
  inv0d0 U8283 ( .I(n8492), .ZN(n3516) );
  nd02d1 U8284 ( .A1(n2988), .A2(n4984), .ZN(n4937) );
  nd02d1 U8285 ( .A1(n9731), .A2(n4974), .ZN(n8227) );
  nd03d1 U8286 ( .A1(n9542), .A2(n2819), .A3(n10359), .ZN(n8792) );
  nd02d1 U8287 ( .A1(N11511), .A2(n5338), .ZN(n7013) );
  inv0d0 U8288 ( .I(n11440), .ZN(n5293) );
  nd02d1 U8289 ( .A1(n12063), .A2(n6871), .ZN(n11493) );
  nr02d1 U8294 ( .A1(n8146), .A2(n4608), .ZN(n9659) );
  nd02d1 U8295 ( .A1(n11534), .A2(n3929), .ZN(n6899) );
  nd02d1 U8298 ( .A1(n11656), .A2(n5259), .ZN(n11661) );
  nd02d1 U8301 ( .A1(N13010), .A2(n12004), .ZN(n9363) );
  nr02d1 U8304 ( .A1(n10262), .A2(n4984), .ZN(n10259) );
  nd02d1 U8305 ( .A1(n4075), .A2(n5203), .ZN(n6799) );
  inv0d0 U8307 ( .I(n8737), .ZN(n3017) );
  inv0d0 U8308 ( .I(n10023), .ZN(n3461) );
  inv0d0 U8309 ( .I(n4955), .ZN(n5729) );
  nd02d1 U8311 ( .A1(n11696), .A2(n3418), .ZN(n4539) );
  nd02d1 U8312 ( .A1(n5829), .A2(n4154), .ZN(n7541) );
  inv0d0 U8313 ( .I(n4772), .ZN(n3098) );
  nd02d1 U8314 ( .A1(n3881), .A2(n10676), .ZN(n7675) );
  nr02d1 U8315 ( .A1(n8430), .A2(n6115), .ZN(n8428) );
  inv0d0 U8317 ( .I(n6106), .ZN(n5544) );
  nd03d1 U8320 ( .A1(n7370), .A2(n3129), .A3(n9453), .ZN(n8669) );
  nd12d1 U8321 ( .A1(n1879), .A2(n11697), .ZN(n8549) );
  inv0d0 U8323 ( .I(n7395), .ZN(n5833) );
  nr02d1 U8324 ( .A1(n5769), .A2(n6935), .ZN(n6627) );
  nr02d1 U8325 ( .A1(n5330), .A2(n7740), .ZN(n7007) );
  nd03d1 U8327 ( .A1(n3076), .A2(n8711), .A3(n3121), .ZN(n8709) );
  nd02d1 U8328 ( .A1(n4086), .A2(n5104), .ZN(n9799) );
  nr02d1 U8331 ( .A1(n4951), .A2(n5757), .ZN(n8421) );
  nd02d1 U8332 ( .A1(n5516), .A2(n4967), .ZN(n5521) );
  nr02d1 U8333 ( .A1(n9931), .A2(n6115), .ZN(n9934) );
  inv0d0 U8334 ( .I(n7955), .ZN(n3116) );
  inv0d0 U8335 ( .I(n5308), .ZN(n4457) );
  nd02d1 U8336 ( .A1(n4442), .A2(n8855), .ZN(n7409) );
  nr02d1 U8337 ( .A1(n3986), .A2(n6650), .ZN(n5954) );
  nd03d1 U8338 ( .A1(n7422), .A2(n8086), .A3(n7420), .ZN(n7676) );
  nd03d1 U8340 ( .A1(n9697), .A2(n5312), .A3(N8380), .ZN(n9700) );
  nr02d1 U8341 ( .A1(n9304), .A2(n8534), .ZN(n7091) );
  inv0d0 U8342 ( .I(n8518), .ZN(n5642) );
  nd02d1 U8343 ( .A1(n4968), .A2(n4639), .ZN(n4644) );
  inv0d0 U8344 ( .I(n4791), .ZN(n3007) );
  nd03d1 U8345 ( .A1(n11182), .A2(n4886), .A3(n2897), .ZN(n8024) );
  inv0d0 U8346 ( .I(n6858), .ZN(n4048) );
  nd02d1 U8347 ( .A1(n3960), .A2(n4958), .ZN(n6930) );
  inv0d0 U8352 ( .I(n10738), .ZN(n3660) );
  inv0d0 U8354 ( .I(n8097), .ZN(n5101) );
  nr02d1 U8356 ( .A1(n6921), .A2(n3961), .ZN(n5178) );
  nr02d1 U8357 ( .A1(n8343), .A2(n5109), .ZN(n6868) );
  inv0d0 U8358 ( .I(n8510), .ZN(n3475) );
  nr02d1 U8359 ( .A1(n10221), .A2(n5231), .ZN(n10223) );
  nr02d1 U8360 ( .A1(n9834), .A2(n5098), .ZN(n9835) );
  inv0d0 U8361 ( .I(n8810), .ZN(n2879) );
  nr02d1 U8362 ( .A1(n8945), .A2(n6070), .ZN(n8946) );
  nr02d1 U8363 ( .A1(n8510), .A2(n5382), .ZN(n7053) );
  nd03d1 U8364 ( .A1(n6421), .A2(n5806), .A3(n3232), .ZN(n7907) );
  nr02d1 U8365 ( .A1(n5576), .A2(n4953), .ZN(n5578) );
  nr02d1 U8366 ( .A1(n6565), .A2(n10819), .ZN(n10830) );
  nr02d1 U8368 ( .A1(n6982), .A2(n5798), .ZN(n7989) );
  nd02d1 U8374 ( .A1(n3418), .A2(n5254), .ZN(n6204) );
  nr02d1 U8375 ( .A1(n6774), .A2(n9775), .ZN(n9779) );
  nr02d1 U8378 ( .A1(n9007), .A2(n6061), .ZN(n9010) );
  nr02d1 U8379 ( .A1(n9855), .A2(n5278), .ZN(n9859) );
  inv0d0 U8382 ( .I(n7447), .ZN(n5458) );
  inv0d0 U8383 ( .I(n11552), .ZN(n3953) );
  nd02d1 U8385 ( .A1(n6319), .A2(n4975), .ZN(n6323) );
  nd02d1 U8386 ( .A1(n7939), .A2(n9471), .ZN(n8692) );
  nd03d1 U8387 ( .A1(n7003), .A2(n7004), .A3(n5544), .ZN(n5323) );
  nd03d1 U8389 ( .A1(n7455), .A2(n8203), .A3(n7456), .ZN(n8207) );
  nr02d1 U8390 ( .A1(n8060), .A2(n4970), .ZN(n7876) );
  inv0d0 U8392 ( .I(n4394), .ZN(n3939) );
  nd02d1 U8393 ( .A1(n8026), .A2(n10326), .ZN(n8027) );
  inv0d0 U8394 ( .I(n7339), .ZN(n2805) );
  inv0d0 U8395 ( .I(n4864), .ZN(n2854) );
  inv0d0 U8396 ( .I(n9525), .ZN(n2993) );
  nd02d1 U8397 ( .A1(n9371), .A2(n3266), .ZN(n9370) );
  nd03d1 U8398 ( .A1(n3556), .A2(n6466), .A3(N12034), .ZN(n6165) );
  nd12d1 U8404 ( .A1(n27), .A2(n8738), .ZN(n8745) );
  nd04d1 U8405 ( .A1(n1342), .A2(n1299), .A3(n1247), .A4(n1569), .ZN(n27) );
  nr02d1 U8406 ( .A1(n6979), .A2(n5797), .ZN(n8018) );
  nr02d1 U8407 ( .A1(n9735), .A2(n6140), .ZN(n9738) );
  nd02d1 U8408 ( .A1(n9232), .A2(n6617), .ZN(n9238) );
  inv0d0 U8409 ( .I(n5600), .ZN(n3120) );
  nd03d1 U8411 ( .A1(n4683), .A2(n7748), .A3(n5743), .ZN(n7755) );
  inv0d0 U8412 ( .I(n4884), .ZN(n2874) );
  nd02d1 U8413 ( .A1(n11680), .A2(n10844), .ZN(n7803) );
  nr02d1 U8414 ( .A1(n6367), .A2(n10118), .ZN(n10392) );
  nr02d1 U8415 ( .A1(n7051), .A2(n5386), .ZN(n7055) );
  nd02d1 U8416 ( .A1(n3942), .A2(n5079), .ZN(n9879) );
  inv0d0 U8417 ( .I(n6896), .ZN(n3927) );
  inv0d0 U8418 ( .I(n5292), .ZN(n3807) );
  inv0d0 U8419 ( .I(n6183), .ZN(n3439) );
  inv0d0 U8421 ( .I(n7090), .ZN(n3458) );
  nd03d1 U8423 ( .A1(n5232), .A2(n5068), .A3(n3875), .ZN(n5236) );
  nr02d1 U8424 ( .A1(n7842), .A2(n8072), .ZN(n7849) );
  inv0d0 U8425 ( .I(n11151), .ZN(n2815) );
  inv0d0 U8426 ( .I(n5112), .ZN(n4962) );
  inv0d0 U8427 ( .I(n9299), .ZN(n4439) );
  nr02d1 U8428 ( .A1(n11244), .A2(n5374), .ZN(n6148) );
  inv0d0 U8429 ( .I(n11225), .ZN(n3167) );
  inv0d0 U8430 ( .I(n4970), .ZN(n3146) );
  nr02d1 U8431 ( .A1(n5521), .A2(n5713), .ZN(n5524) );
  nd02d1 U8432 ( .A1(n7378), .A2(n7210), .ZN(n7220) );
  nd02d1 U8433 ( .A1(n6154), .A2(n8498), .ZN(n4473) );
  inv0d0 U8436 ( .I(n9356), .ZN(n3343) );
  nd02d1 U8437 ( .A1(N12882), .A2(n12007), .ZN(n7137) );
  nd02d1 U8438 ( .A1(n5570), .A2(n7624), .ZN(n7628) );
  nr02d1 U8439 ( .A1(n10187), .A2(n5902), .ZN(n10195) );
  inv0d0 U8441 ( .I(n5948), .ZN(n4006) );
  nd02d1 U8444 ( .A1(n8866), .A2(n8355), .ZN(n8357) );
  nd02d1 U8446 ( .A1(n11517), .A2(n5780), .ZN(n11524) );
  aoim22d1 U8447 ( .A1(n3468), .A2(n5390), .B1(n5391), .B2(n5392), .Z(n5387)
         );
  nd02d1 U8450 ( .A1(n5129), .A2(n4804), .ZN(n9517) );
  inv0d0 U8453 ( .I(n5827), .ZN(n5693) );
  inv0d0 U8454 ( .I(n5209), .ZN(n3845) );
  nd03d1 U8455 ( .A1(n3475), .A2(n6922), .A3(N12130), .ZN(n10013) );
  inv0d0 U8456 ( .I(n8658), .ZN(n3220) );
  inv0d0 U8458 ( .I(n9636), .ZN(n5570) );
  nd03d1 U8459 ( .A1(n3845), .A2(n6861), .A3(N10776), .ZN(n10680) );
  nd03d1 U8461 ( .A1(n4102), .A2(n6547), .A3(n4322), .ZN(n7594) );
  nd02d1 U8464 ( .A1(n6235), .A2(n10893), .ZN(n10897) );
  inv0d0 U8466 ( .I(n10296), .ZN(n2862) );
  inv0d0 U8467 ( .I(n11586), .ZN(n3736) );
  nr02d1 U8468 ( .A1(n11352), .A2(n6884), .ZN(n11355) );
  nd02d1 U8469 ( .A1(n2926), .A2(n11849), .ZN(n4785) );
  inv0d0 U8470 ( .I(n5398), .ZN(n6018) );
  nd02d1 U8471 ( .A1(n3416), .A2(n4663), .ZN(n6210) );
  nd03d1 U8472 ( .A1(n5536), .A2(n4964), .A3(n5711), .ZN(n5561) );
  inv0d0 U8478 ( .I(n5702), .ZN(n5904) );
  inv0d0 U8480 ( .I(n8445), .ZN(n3770) );
  inv0d0 U8482 ( .I(n8312), .ZN(n3996) );
  inv0d0 U8485 ( .I(n7430), .ZN(n5192) );
  nd02d1 U8489 ( .A1(n3456), .A2(n9304), .ZN(n7094) );
  inv0d0 U8490 ( .I(n7998), .ZN(n2914) );
  nd02d1 U8493 ( .A1(n8876), .A2(n11470), .ZN(n7598) );
  nd03d1 U8494 ( .A1(n2863), .A2(n4633), .A3(n11193), .ZN(n9555) );
  inv0d0 U8495 ( .I(n8628), .ZN(n3152) );
  inv0d0 U8496 ( .I(n9606), .ZN(n4305) );
  nr02d1 U8497 ( .A1(n4750), .A2(n4947), .ZN(n4753) );
  nd02d1 U8498 ( .A1(n3832), .A2(n5276), .ZN(n6020) );
  inv0d0 U8500 ( .I(n11196), .ZN(n2984) );
  nd02d1 U8503 ( .A1(n4967), .A2(n3160), .ZN(n4650) );
  inv0d0 U8505 ( .I(n7366), .ZN(n5237) );
  nd02d1 U8506 ( .A1(n8170), .A2(n8126), .ZN(n8172) );
  inv0d0 U8507 ( .I(n5755), .ZN(n5748) );
  nr13d1 U8512 ( .A1(n8884), .A2(n8222), .A3(n8224), .ZN(n8233) );
  inv0d0 U8513 ( .I(n5102), .ZN(n4034) );
  nd02d1 U8517 ( .A1(n9246), .A2(n12040), .ZN(n6137) );
  inv0d0 U8518 ( .I(n7443), .ZN(n5690) );
  inv0d0 U8519 ( .I(n7158), .ZN(n4656) );
  inv0d0 U8520 ( .I(n5917), .ZN(n4078) );
  inv0d0 U8521 ( .I(n5135), .ZN(n3922) );
  inv0d0 U8522 ( .I(n6486), .ZN(n3110) );
  nd02d1 U8523 ( .A1(n5348), .A2(n11250), .ZN(n4395) );
  inv0d0 U8524 ( .I(n7952), .ZN(n3062) );
  inv0d0 U8525 ( .I(n7352), .ZN(n2873) );
  inv0d0 U8526 ( .I(n9990), .ZN(n3507) );
  nd02d1 U8528 ( .A1(n6617), .A2(n4949), .ZN(n7025) );
  inv0d0 U8529 ( .I(n11857), .ZN(n3006) );
  nd02d1 U8530 ( .A1(n3043), .A2(n7923), .ZN(n6578) );
  nd02d1 U8531 ( .A1(n3293), .A2(n5043), .ZN(n6327) );
  inv0d0 U8533 ( .I(n11129), .ZN(n2858) );
  inv0d0 U8534 ( .I(n7845), .ZN(n3251) );
  nd02d1 U8535 ( .A1(n10480), .A2(n6070), .ZN(n9704) );
  inv0d0 U8536 ( .I(n9597), .ZN(n2966) );
  nr13d1 U8537 ( .A1(n4960), .A2(n5709), .A3(n7249), .ZN(n7252) );
  inv0d0 U8538 ( .I(n9953), .ZN(n3774) );
  nd03d1 U8539 ( .A1(n11156), .A2(n5470), .A3(n2885), .ZN(n8009) );
  inv0d0 U8540 ( .I(n9911), .ZN(n3876) );
  nd12d1 U8543 ( .A1(n28), .A2(n6851), .ZN(n6853) );
  aoi21d1 U8544 ( .B1(n1295), .B2(n2358), .A(n1328), .ZN(n28) );
  nd02d1 U8545 ( .A1(n7170), .A2(n7382), .ZN(n7171) );
  inv0d0 U8547 ( .I(n9664), .ZN(n4628) );
  inv0d0 U8549 ( .I(n10368), .ZN(n2967) );
  nd02d1 U8550 ( .A1(n3872), .A2(n6960), .ZN(n9175) );
  inv0d0 U8551 ( .I(n4718), .ZN(n3048) );
  nd02d1 U8552 ( .A1(n3090), .A2(n11973), .ZN(n4761) );
  nd02d1 U8553 ( .A1(n3404), .A2(n4427), .ZN(n6230) );
  nd02d1 U8554 ( .A1(n6808), .A2(n5579), .ZN(n6814) );
  nd03d1 U8555 ( .A1(n3751), .A2(n3761), .A3(n9206), .ZN(n9203) );
  inv0d0 U8556 ( .I(n9212), .ZN(n3712) );
  inv0d0 U8557 ( .I(n10967), .ZN(n3137) );
  nd02d1 U8558 ( .A1(n11993), .A2(n4967), .ZN(n11784) );
  nd02d1 U8559 ( .A1(N12722), .A2(n12015), .ZN(n6217) );
  inv0d0 U8560 ( .I(n1866), .ZN(n1868) );
  nd02d1 U8561 ( .A1(n5362), .A2(n12036), .ZN(n7766) );
  nd02d1 U8562 ( .A1(n3323), .A2(n4653), .ZN(n4585) );
  nd02d1 U8563 ( .A1(n4587), .A2(n5591), .ZN(n10450) );
  nd02d1 U8564 ( .A1(n3962), .A2(n5434), .ZN(n10654) );
  nd02d1 U8565 ( .A1(n4077), .A2(n5957), .ZN(n9062) );
  inv0d0 U8568 ( .I(n9811), .ZN(n4057) );
  nd02d1 U8572 ( .A1(n2836), .A2(n4926), .ZN(n11909) );
  nd02d1 U8573 ( .A1(n2838), .A2(n4926), .ZN(n5686) );
  nd02d1 U8574 ( .A1(n4835), .A2(n6890), .ZN(n11315) );
  nd02d1 U8577 ( .A1(N13522), .A2(n10109), .ZN(n10941) );
  nd02d1 U8578 ( .A1(N12962), .A2(n11726), .ZN(n10892) );
  nd02d1 U8579 ( .A1(n3443), .A2(n4939), .ZN(n7103) );
  nd02d1 U8580 ( .A1(n8554), .A2(n4988), .ZN(n8849) );
  inv0d0 U8581 ( .I(n5289), .ZN(n3748) );
  nd02d1 U8582 ( .A1(N11762), .A2(n12041), .ZN(n10773) );
  nd02d1 U8584 ( .A1(n3312), .A2(n4304), .ZN(n6326) );
  nd02d1 U8585 ( .A1(n11795), .A2(n4964), .ZN(n11797) );
  inv0d0 U8589 ( .I(n10934), .ZN(n3269) );
  inv0d0 U8591 ( .I(n10780), .ZN(n3559) );
  nd02d1 U8592 ( .A1(n2841), .A2(n4926), .ZN(n4867) );
  inv0d0 U8594 ( .I(n11852), .ZN(n3009) );
  inv0d0 U8595 ( .I(n9000), .ZN(n4184) );
  nd02d1 U8596 ( .A1(n4844), .A2(n5714), .ZN(n8132) );
  nd02d1 U8597 ( .A1(N12738), .A2(n11710), .ZN(n9333) );
  inv0d0 U8603 ( .I(n1863), .ZN(n1865) );
  nd02d1 U8604 ( .A1(n10403), .A2(n5348), .ZN(n8465) );
  inv0d0 U8605 ( .I(n4975), .ZN(n5520) );
  inv0d0 U8608 ( .I(n11159), .ZN(n2908) );
  nd02d1 U8609 ( .A1(N12610), .A2(n5422), .ZN(n10049) );
  inv0d0 U8610 ( .I(n9677), .ZN(n4352) );
  inv0d0 U8613 ( .I(n9790), .ZN(n4060) );
  nd02d1 U8614 ( .A1(n8168), .A2(n4368), .ZN(n7486) );
  nd02d1 U8615 ( .A1(n8900), .A2(n6072), .ZN(n9656) );
  inv0d0 U8616 ( .I(n5139), .ZN(n6045) );
  nd02d1 U8618 ( .A1(N12626), .A2(n10054), .ZN(n10057) );
  inv0d0 U8619 ( .I(n1882), .ZN(N12626) );
  inv0d0 U8620 ( .I(n1880), .ZN(n1883) );
  nd02d1 U8621 ( .A1(n3933), .A2(n4464), .ZN(n5151) );
  nd02d1 U8622 ( .A1(n5157), .A2(n3933), .ZN(n5993) );
  nd02d1 U8623 ( .A1(n8075), .A2(n9616), .ZN(n9279) );
  nd02d1 U8624 ( .A1(n3302), .A2(n5370), .ZN(n7198) );
  inv0d0 U8625 ( .I(n11984), .ZN(n3195) );
  inv0d0 U8626 ( .I(n8654), .ZN(n3151) );
  inv0d0 U8627 ( .I(n6604), .ZN(n5406) );
  nd02d1 U8629 ( .A1(n8417), .A2(n5431), .ZN(n11257) );
  inv0d0 U8632 ( .I(n11955), .ZN(n2896) );
  buffd1 U8633 ( .I(n1036), .Z(n1034) );
  inv0d0 U8637 ( .I(n10492), .ZN(n4295) );
  nd02d1 U8638 ( .A1(n3449), .A2(n5405), .ZN(n7102) );
  inv0d0 U8640 ( .I(n11980), .ZN(n3050) );
  inv0d0 U8643 ( .I(n6631), .ZN(n5435) );
  nd02d1 U8644 ( .A1(n3566), .A2(n5168), .ZN(n8477) );
  inv0d0 U8646 ( .I(n10041), .ZN(n3482) );
  inv0d0 U8647 ( .I(n6966), .ZN(n3810) );
  inv0d0 U8649 ( .I(n5330), .ZN(n5837) );
  inv0d0 U8651 ( .I(n9578), .ZN(n2889) );
  nd02d1 U8652 ( .A1(N9470), .A2(n10568), .ZN(n5930) );
  inv0d0 U8654 ( .I(n7085), .ZN(n3436) );
  inv0d0 U8656 ( .I(n10592), .ZN(n3988) );
  nd03d1 U8661 ( .A1(n11955), .A2(n5320), .A3(n11175), .ZN(n8823) );
  inv0d0 U8662 ( .I(n10823), .ZN(n3466) );
  inv0d0 U8665 ( .I(n11371), .ZN(n4330) );
  inv0d0 U8666 ( .I(n11212), .ZN(n3020) );
  inv0d0 U8667 ( .I(n6935), .ZN(n3821) );
  inv0d0 U8668 ( .I(n7583), .ZN(n4083) );
  inv0d0 U8675 ( .I(n11584), .ZN(n3618) );
  inv0d0 U8677 ( .I(n7452), .ZN(n4205) );
  inv0d0 U8678 ( .I(n10086), .ZN(n3272) );
  inv0d0 U8684 ( .I(n10452), .ZN(n4590) );
  aoim22d1 U8686 ( .A1(n7331), .A2(n4933), .B1(n11967), .B2(n4840), .Z(n4848)
         );
  nr02d1 U8689 ( .A1(n11196), .A2(n11966), .ZN(n11967) );
  inv0d0 U8691 ( .I(n6554), .ZN(n5344) );
  nr02d1 U8692 ( .A1(n5005), .A2(n12038), .ZN(n11639) );
  inv0d0 U8693 ( .I(n11062), .ZN(n3104) );
  inv0d0 U8696 ( .I(n10711), .ZN(n3664) );
  inv0d0 U8697 ( .I(n9496), .ZN(n3013) );
  inv0d0 U8702 ( .I(n8694), .ZN(n5621) );
  inv0d0 U8703 ( .I(n5726), .ZN(n5634) );
  nd02d1 U8704 ( .A1(n9425), .A2(n5625), .ZN(n8627) );
  nd02d1 U8705 ( .A1(N14226), .A2(n9459), .ZN(n9461) );
  inv0d0 U8706 ( .I(n9999), .ZN(n3506) );
  nd02d1 U8707 ( .A1(n9586), .A2(n10298), .ZN(n10300) );
  nd02d1 U8709 ( .A1(n8581), .A2(n10086), .ZN(n9374) );
  inv0d0 U8710 ( .I(n7429), .ZN(n4470) );
  inv0d0 U8714 ( .I(n5048), .ZN(n4055) );
  inv0d0 U8719 ( .I(n7382), .ZN(n5631) );
  inv0d0 U8725 ( .I(n4969), .ZN(n4913) );
  nd02d1 U8728 ( .A1(n8862), .A2(n9921), .ZN(n9923) );
  inv0d0 U8732 ( .I(n8424), .ZN(n3864) );
  inv0d0 U8733 ( .I(n8970), .ZN(n4284) );
  inv0d0 U8736 ( .I(n9193), .ZN(n3719) );
  inv0d0 U8740 ( .I(n11973), .ZN(n3112) );
  nd02d1 U8742 ( .A1(n11417), .A2(n7554), .ZN(n11415) );
  inv0d0 U8743 ( .I(n9477), .ZN(n3115) );
  inv0d0 U8744 ( .I(n11268), .ZN(n3904) );
  nd02d1 U8745 ( .A1(n4964), .A2(n4669), .ZN(n4670) );
  inv0d0 U8746 ( .I(n11279), .ZN(n4121) );
  nd02d1 U8747 ( .A1(n3684), .A2(n6617), .ZN(n6124) );
  inv0d0 U8748 ( .I(n8858), .ZN(n5182) );
  inv0d0 U8749 ( .I(n10535), .ZN(n4140) );
  inv0d0 U8750 ( .I(n8933), .ZN(n4346) );
  inv0d0 U8751 ( .I(n7547), .ZN(n4207) );
  nr02d1 U8752 ( .A1(n8688), .A2(n6599), .ZN(n11016) );
  inv0d0 U8753 ( .I(n6034), .ZN(n3839) );
  inv0d0 U8754 ( .I(n6415), .ZN(n4303) );
  inv0d0 U8755 ( .I(n5956), .ZN(n3997) );
  nr02d1 U8756 ( .A1(n8787), .A2(n10276), .ZN(n10275) );
  inv0d0 U8757 ( .I(n6608), .ZN(n4677) );
  inv0d0 U8758 ( .I(n10509), .ZN(n4293) );
  nd03d1 U8759 ( .A1(n11039), .A2(n4406), .A3(n3074), .ZN(n5593) );
  inv0d0 U8762 ( .I(n8109), .ZN(n4323) );
  inv0d0 U8763 ( .I(n11266), .ZN(n3905) );
  inv0d0 U8765 ( .I(n11838), .ZN(n3114) );
  nd02d1 U8766 ( .A1(n6651), .A2(n8302), .ZN(n8304) );
  nd02d1 U8777 ( .A1(n6651), .A2(n5941), .ZN(n5946) );
  inv0d0 U8781 ( .I(n5513), .ZN(n3247) );
  inv0d0 U8783 ( .I(n11143), .ZN(n2816) );
  nd03d1 U8784 ( .A1(n3005), .A2(n10226), .A3(n2944), .ZN(n10225) );
  inv0d0 U8785 ( .I(n9511), .ZN(n2949) );
  nr13d1 U8787 ( .A1(n8857), .A2(n5835), .A3(n9219), .ZN(n9226) );
  inv0d0 U8788 ( .I(n5700), .ZN(n4301) );
  inv0d0 U8789 ( .I(n10361), .ZN(n2973) );
  nd02d1 U8790 ( .A1(n3401), .A2(n8563), .ZN(n6231) );
  inv0d0 U8791 ( .I(n6318), .ZN(n4421) );
  inv0d0 U8792 ( .I(n7517), .ZN(n4257) );
  inv0d0 U8794 ( .I(n8937), .ZN(n4239) );
  nd02d1 U8796 ( .A1(n3343), .A2(n5723), .ZN(n9361) );
  nd02d1 U8797 ( .A1(n5213), .A2(n9706), .ZN(n9708) );
  inv0d0 U8798 ( .I(n9847), .ZN(n4039) );
  nd02d1 U8799 ( .A1(n8161), .A2(n5466), .ZN(n7484) );
  inv0d0 U8800 ( .I(n7896), .ZN(n3156) );
  inv0d0 U8801 ( .I(n8159), .ZN(n4392) );
  inv0d0 U8803 ( .I(n6955), .ZN(n3846) );
  nr02d1 U8805 ( .A1(n10934), .A2(n6293), .ZN(n10933) );
  inv0d0 U8806 ( .I(n8434), .ZN(n3675) );
  inv0d0 U8809 ( .I(n6095), .ZN(n3775) );
  inv0d0 U8811 ( .I(n7350), .ZN(n2853) );
  aoim22d1 U8812 ( .A1(n4103), .A2(n6807), .B1(n5923), .B2(n6808), .Z(n6804)
         );
  inv0d0 U8814 ( .I(n5026), .ZN(n4103) );
  inv0d0 U8815 ( .I(n8121), .ZN(n4291) );
  inv0d0 U8816 ( .I(n7396), .ZN(n4308) );
  inv0d0 U8817 ( .I(n5754), .ZN(n5274) );
  inv0d0 U8818 ( .I(n9903), .ZN(n3835) );
  inv0d0 U8819 ( .I(n11503), .ZN(n4052) );
  inv0d0 U8820 ( .I(n7692), .ZN(n3888) );
  inv0d0 U8822 ( .I(n4591), .ZN(n5252) );
  inv0d0 U8823 ( .I(n9015), .ZN(n4142) );
  inv0d0 U8824 ( .I(n8951), .ZN(n4285) );
  inv0d0 U8825 ( .I(n11891), .ZN(n2825) );
  inv0d0 U8826 ( .I(n4526), .ZN(n3345) );
  inv0d0 U8827 ( .I(n5342), .ZN(n3791) );
  inv0d0 U8828 ( .I(n11187), .ZN(n2882) );
  nr13d1 U8829 ( .A1(n7450), .A2(n5581), .A3(n6755), .ZN(n6760) );
  inv0d0 U8830 ( .I(n7762), .ZN(n3561) );
  nr13d1 U8831 ( .A1(n7317), .A2(n7314), .A3(n5126), .ZN(n7320) );
  inv0d0 U8832 ( .I(n5936), .ZN(n4322) );
  inv0d0 U8833 ( .I(n10843), .ZN(n3485) );
  inv0d0 U8834 ( .I(n8606), .ZN(n3305) );
  inv0d0 U8835 ( .I(n6313), .ZN(n3283) );
  inv0d0 U8836 ( .I(n6680), .ZN(n5794) );
  inv0d0 U8837 ( .I(n5859), .ZN(n4172) );
  inv0d0 U8838 ( .I(n8162), .ZN(n4339) );
  inv0d0 U8839 ( .I(n11158), .ZN(n2814) );
  nd02d1 U8840 ( .A1(n4154), .A2(n5204), .ZN(n8249) );
  nd02d1 U8841 ( .A1(n8633), .A2(n4964), .ZN(n8643) );
  inv0d0 U8842 ( .I(n8014), .ZN(n2890) );
  inv0d0 U8843 ( .I(n6733), .ZN(n4216) );
  inv0d0 U8844 ( .I(n10850), .ZN(n3421) );
  inv0d0 U8845 ( .I(n6014), .ZN(n3826) );
  nd02d1 U8846 ( .A1(n5465), .A2(n8220), .ZN(n8224) );
  inv0d0 U8847 ( .I(n4611), .ZN(n5152) );
  nd02d1 U8848 ( .A1(n6783), .A2(n4116), .ZN(n5885) );
  inv0d0 U8849 ( .I(n5967), .ZN(n4025) );
  inv0d0 U8850 ( .I(n11828), .ZN(n3061) );
  nr13d1 U8851 ( .A1(n5720), .A2(n3260), .A3(n6294), .ZN(n8591) );
  inv0d0 U8852 ( .I(n5234), .ZN(n5550) );
  inv0d0 U8853 ( .I(n5905), .ZN(n4111) );
  inv0d0 U8854 ( .I(n9259), .ZN(n3558) );
  nr02d1 U8855 ( .A1(n10379), .A2(n3118), .ZN(n10196) );
  inv0d0 U8856 ( .I(n8712), .ZN(n3118) );
  inv0d0 U8857 ( .I(n8828), .ZN(n2911) );
  inv0d0 U8858 ( .I(n11835), .ZN(n3080) );
  inv0d0 U8859 ( .I(n4982), .ZN(n4922) );
  inv0d0 U8860 ( .I(n6421), .ZN(n3233) );
  inv0d0 U8862 ( .I(n10504), .ZN(n4294) );
  inv0d0 U8863 ( .I(n4924), .ZN(n5124) );
  inv0d0 U8864 ( .I(n7436), .ZN(n5687) );
  inv0d0 U8865 ( .I(n9640), .ZN(n3991) );
  nr13d1 U8866 ( .A1(n4956), .A2(n6160), .A3(n6429), .ZN(n6574) );
  nd02d1 U8868 ( .A1(n3936), .A2(n5558), .ZN(n7659) );
  nd02d1 U8869 ( .A1(n5705), .A2(n6890), .ZN(n8139) );
  nd02d1 U8870 ( .A1(n11637), .A2(n6618), .ZN(n9240) );
  nd02d1 U8871 ( .A1(n3969), .A2(n9848), .ZN(n5984) );
  inv0d0 U8872 ( .I(n4993), .ZN(n4941) );
  nr13d1 U8873 ( .A1(n5724), .A2(n6297), .A3(n5446), .ZN(n5452) );
  inv0d0 U8874 ( .I(n8813), .ZN(n2886) );
  nr13d1 U8875 ( .A1(n7388), .A2(n4982), .A3(n7140), .ZN(n7145) );
  inv0d0 U8876 ( .I(n6823), .ZN(n4093) );
  inv0d0 U8877 ( .I(n9679), .ZN(n4357) );
  inv0d0 U8878 ( .I(n10455), .ZN(n4549) );
  inv0d0 U8879 ( .I(n11259), .ZN(n3878) );
  inv0d0 U8880 ( .I(n8475), .ZN(n5647) );
  nd02d1 U8881 ( .A1(n3298), .A2(n4902), .ZN(n8843) );
  nd02d1 U8883 ( .A1(n5734), .A2(n9612), .ZN(n9328) );
  inv0d0 U8884 ( .I(n7578), .ZN(n4075) );
  inv0d0 U8885 ( .I(n7413), .ZN(n5655) );
  inv0d0 U8886 ( .I(n6417), .ZN(n3234) );
  inv0d0 U8888 ( .I(n8473), .ZN(n3533) );
  inv0d0 U8890 ( .I(n6713), .ZN(n4250) );
  inv0d0 U8891 ( .I(n8074), .ZN(n5734) );
  inv0d0 U8892 ( .I(n10319), .ZN(n2824) );
  inv0d0 U8893 ( .I(n10326), .ZN(n2904) );
  inv0d0 U8894 ( .I(n10445), .ZN(n4819) );
  inv0d0 U8895 ( .I(n6402), .ZN(n5518) );
  inv0d0 U8896 ( .I(n10632), .ZN(n3965) );
  inv0d0 U8898 ( .I(n5866), .ZN(n4167) );
  inv0d0 U8899 ( .I(n5430), .ZN(n3338) );
  inv0d0 U8900 ( .I(n4660), .ZN(n3182) );
  inv0d0 U8902 ( .I(n10045), .ZN(n3445) );
  inv0d0 U8907 ( .I(n12052), .ZN(n3866) );
  inv0d0 U8909 ( .I(n9197), .ZN(n4693) );
  inv0d0 U8911 ( .I(n10630), .ZN(n3921) );
  inv0d0 U8912 ( .I(n5961), .ZN(n4056) );
  inv0d0 U8913 ( .I(n8214), .ZN(n4259) );
  buffd1 U8914 ( .I(n1086), .Z(n1043) );
  inv0d0 U8915 ( .I(n5193), .ZN(n3817) );
  buffd1 U8918 ( .I(n1086), .Z(n1042) );
  inv0d0 U8919 ( .I(n5109), .ZN(n4044) );
  inv0d0 U8920 ( .I(n5981), .ZN(n3968) );
  nd02d1 U8921 ( .A1(n11572), .A2(n6624), .ZN(n11576) );
  inv0d0 U8922 ( .I(n10486), .ZN(n4276) );
  inv0d0 U8923 ( .I(n4953), .ZN(n4646) );
  inv0d0 U8924 ( .I(n4963), .ZN(n5910) );
  nd02d1 U8926 ( .A1(n8611), .A2(n4913), .ZN(n8834) );
  inv0d0 U8927 ( .I(n10931), .ZN(n3289) );
  inv0d0 U8928 ( .I(n5296), .ZN(n6033) );
  inv0d0 U8929 ( .I(n9574), .ZN(n2892) );
  inv0d0 U8930 ( .I(n7028), .ZN(n3566) );
  inv0d0 U8931 ( .I(n8752), .ZN(n2957) );
  inv0d0 U8932 ( .I(n7427), .ZN(n5096) );
  inv0d0 U8933 ( .I(n12043), .ZN(n3528) );
  inv0d0 U8934 ( .I(n9050), .ZN(n4066) );
  inv0d0 U8936 ( .I(n5218), .ZN(n4462) );
  inv0d0 U8937 ( .I(n5742), .ZN(n5061) );
  inv0d0 U8938 ( .I(n5757), .ZN(n5433) );
  inv0d0 U8939 ( .I(n9542), .ZN(n2831) );
  inv0d0 U8941 ( .I(n10020), .ZN(n3470) );
  inv0d0 U8942 ( .I(n6619), .ZN(n5939) );
  inv0d0 U8943 ( .I(n8033), .ZN(n2934) );
  inv0d0 U8945 ( .I(n8874), .ZN(n4095) );
  nd02d1 U8946 ( .A1(n4966), .A2(n6834), .ZN(n8875) );
  inv0d0 U8947 ( .I(n11378), .ZN(n4266) );
  inv0d0 U8948 ( .I(n5246), .ZN(n3854) );
  inv0d0 U8949 ( .I(n6789), .ZN(n4070) );
  inv0d0 U8950 ( .I(n11689), .ZN(n3362) );
  inv0d0 U8951 ( .I(n7131), .ZN(n3353) );
  inv0d0 U8953 ( .I(n11022), .ZN(n3126) );
  inv0d0 U8955 ( .I(n7599), .ZN(n4092) );
  inv0d0 U8956 ( .I(n4990), .ZN(n4668) );
  inv0d0 U8957 ( .I(n10428), .ZN(n4619) );
  inv0d0 U8959 ( .I(n8704), .ZN(n3077) );
  inv0d0 U8960 ( .I(n5121), .ZN(n3967) );
  inv0d0 U8962 ( .I(n10004), .ZN(n3484) );
  inv0d0 U8963 ( .I(n8082), .ZN(n4954) );
  inv0d0 U8964 ( .I(n6649), .ZN(n3995) );
  buffd1 U8965 ( .I(n997), .Z(n984) );
  inv0d0 U8966 ( .I(n957), .ZN(n997) );
  inv0d0 U8967 ( .I(n8863), .ZN(n5071) );
  inv0d0 U8968 ( .I(n6825), .ZN(n5449) );
  inv0d0 U8969 ( .I(n9638), .ZN(n4008) );
  inv0d0 U8970 ( .I(n5803), .ZN(n5779) );
  inv0d0 U8971 ( .I(n5713), .ZN(n5987) );
  inv0d0 U8972 ( .I(n10984), .ZN(n3186) );
  inv0d0 U8973 ( .I(n8251), .ZN(n4156) );
  inv0d0 U8975 ( .I(n8323), .ZN(n4022) );
  inv0d0 U8976 ( .I(n7434), .ZN(n5441) );
  inv0d0 U8978 ( .I(n9471), .ZN(n3125) );
  inv0d0 U8980 ( .I(n6696), .ZN(n4275) );
  inv0d0 U8981 ( .I(n5481), .ZN(n3253) );
  inv0d0 U8982 ( .I(n8093), .ZN(n4711) );
  inv0d0 U8983 ( .I(n6874), .ZN(n3966) );
  inv0d0 U8984 ( .I(n6296), .ZN(n5997) );
  inv0d0 U8985 ( .I(n10932), .ZN(n3288) );
  inv0d0 U8986 ( .I(n8759), .ZN(n5129) );
  inv0d0 U8987 ( .I(n7376), .ZN(n3196) );
  inv0d0 U8988 ( .I(n6394), .ZN(n3200) );
  inv0d0 U8989 ( .I(n7481), .ZN(n5870) );
  inv0d0 U8990 ( .I(n11434), .ZN(n4115) );
  inv0d0 U8991 ( .I(n8977), .ZN(n5465) );
  inv0d0 U8992 ( .I(n8373), .ZN(n3944) );
  inv0d0 U8993 ( .I(n11903), .ZN(n6079) );
  inv0d0 U8994 ( .I(n7704), .ZN(n4315) );
  inv0d0 U8995 ( .I(n5144), .ZN(n3924) );
  inv0d0 U8996 ( .I(n7502), .ZN(n4273) );
  inv0d0 U8997 ( .I(n8290), .ZN(n4080) );
  inv0d0 U8998 ( .I(n7457), .ZN(n5213) );
  inv0d0 U8999 ( .I(n7918), .ZN(n3044) );
  inv0d0 U9000 ( .I(n6594), .ZN(n3161) );
  inv0d0 U9001 ( .I(n8979), .ZN(n4268) );
  inv0d0 U9003 ( .I(n11390), .ZN(n4199) );
  inv0d0 U9004 ( .I(n10243), .ZN(n2918) );
  inv0d0 U9005 ( .I(n5741), .ZN(n4309) );
  inv0d0 U9007 ( .I(n11997), .ZN(n3246) );
  inv0d0 U9008 ( .I(n6662), .ZN(n5582) );
  inv0d0 U9010 ( .I(n5256), .ZN(n3861) );
  inv0d0 U9011 ( .I(n5454), .ZN(n3336) );
  inv0d0 U9012 ( .I(n7433), .ZN(n5683) );
  inv0d0 U9013 ( .I(n6612), .ZN(n5413) );
  inv0d0 U9014 ( .I(n6885), .ZN(n4719) );
  inv0d0 U9015 ( .I(n10416), .ZN(n4742) );
  inv0d0 U9016 ( .I(n5358), .ZN(n3540) );
  inv0d0 U9017 ( .I(n12033), .ZN(n5414) );
  inv0d0 U9018 ( .I(n5769), .ZN(n4957) );
  inv0d0 U9020 ( .I(n5054), .ZN(n5771) );
  inv0d0 U9021 ( .I(n11325), .ZN(n4572) );
  inv0d0 U9022 ( .I(n4947), .ZN(n5495) );
  inv0d0 U9023 ( .I(n8781), .ZN(n2977) );
  inv0d0 U9026 ( .I(n7400), .ZN(n5052) );
  inv0d0 U9027 ( .I(n10230), .ZN(n2951) );
  inv0d0 U9028 ( .I(n7149), .ZN(n3327) );
  inv0d0 U9029 ( .I(n11244), .ZN(n3548) );
  inv0d0 U9030 ( .I(n4997), .ZN(n3426) );
  inv0d0 U9031 ( .I(n11860), .ZN(n2950) );
  inv0d0 U9032 ( .I(n7375), .ZN(n5035) );
  inv0d0 U9033 ( .I(n8370), .ZN(n5567) );
  inv0d0 U9034 ( .I(n7585), .ZN(n4106) );
  aoim22d1 U9035 ( .A1(n3536), .A2(n8484), .B1(n12040), .B2(n3564), .Z(n9248)
         );
  inv0d0 U9036 ( .I(n8992), .ZN(n4224) );
  inv0d0 U9037 ( .I(n7640), .ZN(n5442) );
  inv0d0 U9038 ( .I(n5167), .ZN(n3938) );
  inv0d0 U9039 ( .I(n9691), .ZN(n4296) );
  aoim22d1 U9040 ( .A1(n6591), .A2(n8634), .B1(n8635), .B2(n3183), .Z(n4661)
         );
  inv0d0 U9041 ( .I(n6774), .ZN(n6139) );
  inv0d0 U9042 ( .I(n6611), .ZN(n3503) );
  inv0d0 U9044 ( .I(n12030), .ZN(n3546) );
  inv0d0 U9045 ( .I(n6685), .ZN(n5784) );
  inv0d0 U9046 ( .I(n5386), .ZN(n5259) );
  aoim22d1 U9047 ( .A1(n9437), .A2(n5506), .B1(n11803), .B2(n11804), .Z(n7899)
         );
  nd02d1 U9048 ( .A1(n3206), .A2(n5034), .ZN(n11804) );
  inv0d0 U9049 ( .I(n9628), .ZN(n3892) );
  inv0d0 U9050 ( .I(n10459), .ZN(n4561) );
  inv0d0 U9054 ( .I(n5332), .ZN(n3783) );
  inv0d0 U9055 ( .I(n8311), .ZN(n4003) );
  inv0d0 U9056 ( .I(n7209), .ZN(n3169) );
  inv0d0 U9057 ( .I(n9011), .ZN(n5697) );
  inv0d0 U9058 ( .I(n8463), .ZN(n3571) );
  inv0d0 U9059 ( .I(n6399), .ZN(n3142) );
  inv0d0 U9060 ( .I(n5733), .ZN(n4437) );
  inv0d0 U9062 ( .I(n6622), .ZN(n6117) );
  inv0d0 U9063 ( .I(n7619), .ZN(n4020) );
  inv0d0 U9064 ( .I(n5816), .ZN(n4183) );
  inv0d0 U9065 ( .I(n8275), .ZN(n4128) );
  inv0d0 U9066 ( .I(n11613), .ZN(n3778) );
  inv0d0 U9067 ( .I(n11194), .ZN(n2859) );
  inv0d0 U9068 ( .I(n5099), .ZN(n4037) );
  inv0d0 U9070 ( .I(n11253), .ZN(n3527) );
  inv0d0 U9071 ( .I(n8020), .ZN(n4889) );
  inv0d0 U9072 ( .I(n8129), .ZN(n4767) );
  inv0d0 U9073 ( .I(n11561), .ZN(n5756) );
  inv0d0 U9074 ( .I(n10363), .ZN(n2916) );
  inv0d0 U9075 ( .I(n8815), .ZN(n4396) );
  inv0d0 U9076 ( .I(n6921), .ZN(n5849) );
  buffd1 U9077 ( .I(n1372), .Z(n1368) );
  buffd1 U9078 ( .I(n1372), .Z(n1369) );
  buffd1 U9079 ( .I(n1039), .Z(n1080) );
  buffd1 U9080 ( .I(n1372), .Z(n1366) );
  buffd1 U9081 ( .I(n1372), .Z(n1370) );
  buffd1 U9082 ( .I(n1372), .Z(n1371) );
  buffd1 U9083 ( .I(n1372), .Z(n1367) );
  buffd1 U9084 ( .I(n1040), .Z(n1084) );
  buffd1 U9085 ( .I(n1039), .Z(n1082) );
  buffd1 U9086 ( .I(n1038), .Z(n1078) );
  buffd1 U9087 ( .I(n1040), .Z(n1083) );
  buffd1 U9088 ( .I(n1038), .Z(n1077) );
  buffd1 U9089 ( .I(n1037), .Z(n1076) );
  buffd1 U9090 ( .I(n1040), .Z(n1085) );
  buffd1 U9091 ( .I(n1039), .Z(n1081) );
  buffd1 U9092 ( .I(n1037), .Z(n1075) );
  buffd1 U9093 ( .I(n1037), .Z(n1074) );
  buffd1 U9094 ( .I(n1038), .Z(n1079) );
  buffd1 U9096 ( .I(n7567), .Z(n546) );
  buffd1 U9097 ( .I(n7567), .Z(n549) );
  buffd1 U9098 ( .I(n7567), .Z(n547) );
  buffd1 U9099 ( .I(n7567), .Z(n548) );
  buffd1 U9100 ( .I(n707), .Z(n659) );
  buffd1 U9101 ( .I(n550), .Z(n707) );
  buffd1 U9102 ( .I(n7567), .Z(n550) );
  inv0d0 U9104 ( .I(n7974), .ZN(n4895) );
  inv0d0 U9105 ( .I(n8767), .ZN(n4405) );
  inv0d0 U9106 ( .I(n10430), .ZN(n4827) );
  inv0d0 U9107 ( .I(n5774), .ZN(n4317) );
  inv0d0 U9108 ( .I(n5786), .ZN(n4471) );
  inv0d0 U9110 ( .I(n10587), .ZN(n4000) );
  inv0d0 U9111 ( .I(n11571), .ZN(n3838) );
  inv0d0 U9112 ( .I(n9657), .ZN(n4847) );
  inv0d0 U9113 ( .I(n8903), .ZN(n5705) );
  inv0d0 U9114 ( .I(n8575), .ZN(n3392) );
  inv0d0 U9115 ( .I(n8250), .ZN(n4219) );
  inv0d0 U9116 ( .I(n10453), .ZN(n4595) );
  buffd1 U9117 ( .I(n1036), .Z(n1035) );
  inv0d0 U9118 ( .I(n4519), .ZN(n3500) );
  inv0d0 U9119 ( .I(n10210), .ZN(n3134) );
  inv0d0 U9120 ( .I(n5421), .ZN(n3480) );
  inv0d0 U9121 ( .I(n7473), .ZN(n5595) );
  inv0d0 U9122 ( .I(n8111), .ZN(n4209) );
  inv0d0 U9123 ( .I(n9625), .ZN(n5652) );
  inv0d0 U9124 ( .I(n8901), .ZN(n4866) );
  inv0d0 U9125 ( .I(n10347), .ZN(n2822) );
  inv0d0 U9126 ( .I(n9123), .ZN(n3981) );
  inv0d0 U9127 ( .I(n7368), .ZN(n3221) );
  inv0d0 U9128 ( .I(n11311), .ZN(n4844) );
  inv0d0 U9129 ( .I(n6468), .ZN(n4408) );
  inv0d0 U9130 ( .I(n11880), .ZN(n4299) );
  inv0d0 U9131 ( .I(n8512), .ZN(n5165) );
  inv0d0 U9132 ( .I(n11451), .ZN(n2790) );
  inv0d0 U9133 ( .I(n10413), .ZN(n5763) );
  inv0d0 U9134 ( .I(n10412), .ZN(n4725) );
  inv0d0 U9135 ( .I(n9338), .ZN(n3344) );
  aoim22d1 U9136 ( .A1(n7997), .A2(n7998), .B1(n7999), .B2(n2829), .Z(n7996)
         );
  inv0d0 U9137 ( .I(n10397), .ZN(n4312) );
  nr13d1 U9139 ( .A1(n5511), .A2(n5513), .A3(n5514), .ZN(n5509) );
  aoim22d1 U9140 ( .A1(n2905), .A2(n6508), .B1(n4891), .B2(n4297), .Z(n9572)
         );
  inv0d0 U9141 ( .I(n5439), .ZN(n3337) );
  inv0d0 U9142 ( .I(n9341), .ZN(n3341) );
  inv0d0 U9143 ( .I(n8560), .ZN(n2795) );
  inv0d0 U9144 ( .I(n5766), .ZN(n5753) );
  inv0d0 U9145 ( .I(n8878), .ZN(n4126) );
  inv0d0 U9146 ( .I(n9681), .ZN(n4347) );
  inv0d0 U9147 ( .I(n9054), .ZN(n4137) );
  inv0d0 U9148 ( .I(n10351), .ZN(n2821) );
  inv0d0 U9149 ( .I(n9405), .ZN(n3262) );
  inv0d0 U9151 ( .I(n7051), .ZN(n3486) );
  inv0d0 U9152 ( .I(n9163), .ZN(n3893) );
  inv0d0 U9153 ( .I(n6298), .ZN(n3276) );
  inv0d0 U9154 ( .I(n1270), .ZN(n1321) );
  inv0d0 U9155 ( .I(n1270), .ZN(n1320) );
  inv0d0 U9156 ( .I(n1221), .ZN(n1268) );
  inv0d0 U9157 ( .I(n957), .ZN(n995) );
  inv0d0 U9159 ( .I(n1221), .ZN(n1267) );
  inv0d0 U9160 ( .I(n1270), .ZN(n1322) );
  inv0d0 U9161 ( .I(n957), .ZN(n996) );
  inv0d0 U9162 ( .I(n1221), .ZN(n1266) );
  inv0d0 U9163 ( .I(n957), .ZN(n994) );
  inv0d0 U9164 ( .I(n1132), .ZN(n1174) );
  inv0d0 U9165 ( .I(n1175), .ZN(n1218) );
  inv0d0 U9166 ( .I(n1132), .ZN(n1172) );
  inv0d0 U9168 ( .I(n1175), .ZN(n1219) );
  inv0d0 U9169 ( .I(n1175), .ZN(n1220) );
  inv0d0 U9170 ( .I(n1132), .ZN(n1173) );
  inv0d0 U9171 ( .I(n1087), .ZN(n1129) );
  inv0d0 U9175 ( .I(n1087), .ZN(n1130) );
  inv0d0 U9176 ( .I(n10064), .ZN(n3332) );
  inv0d0 U9177 ( .I(n9801), .ZN(n4058) );
  inv0d0 U9178 ( .I(n1270), .ZN(n1323) );
  inv0d0 U9179 ( .I(n1087), .ZN(n1131) );
  inv0d1 U9181 ( .I(reorder_O2[4]), .ZN(n7293) );
  inv0d1 U9182 ( .I(reorder_O2[1]), .ZN(n7377) );
  inv0d1 U9183 ( .I(reorder_O2[5]), .ZN(n7288) );
  inv0d1 U9184 ( .I(reorder_O2[6]), .ZN(n7278) );
  inv0d1 U9185 ( .I(reorder_O2[0]), .ZN(n7408) );
  inv0d1 U9186 ( .I(reorder_O2[2]), .ZN(n7318) );
  inv0d1 U9187 ( .I(reorder_O2[3]), .ZN(n7297) );
  inv0d1 U9188 ( .I(reorder_O2[7]), .ZN(n7271) );
  inv0d1 U9189 ( .I(reorder_O2[10]), .ZN(n7405) );
  inv0d1 U9190 ( .I(reorder_O2[9]), .ZN(n7261) );
  inv0d1 U9192 ( .I(reorder_O2[20]), .ZN(n7372) );
  inv0d1 U9193 ( .I(reorder_O2[30]), .ZN(n7312) );
  inv0d1 U9194 ( .I(reorder_O2[14]), .ZN(n7398) );
  inv0d1 U9195 ( .I(reorder_O2[21]), .ZN(n7371) );
  inv0d1 U9196 ( .I(reorder_O2[24]), .ZN(n7361) );
  inv0d1 U9197 ( .I(reorder_O2[27]), .ZN(n7342) );
  inv0d1 U9198 ( .I(reorder_O2[8]), .ZN(n7265) );
  inv0d1 U9199 ( .I(reorder_O2[11]), .ZN(n7403) );
  inv0d1 U9200 ( .I(reorder_O2[19]), .ZN(n7379) );
  inv0d1 U9201 ( .I(reorder_O2[12]), .ZN(n7402) );
  inv0d1 U9202 ( .I(reorder_O2[13]), .ZN(n7399) );
  inv0d1 U9203 ( .I(reorder_O2[15]), .ZN(n7397) );
  inv0d1 U9204 ( .I(reorder_O2[16]), .ZN(n7390) );
  inv0d1 U9205 ( .I(reorder_O2[17]), .ZN(n7387) );
  inv0d1 U9206 ( .I(reorder_O2[18]), .ZN(n7380) );
  inv0d1 U9207 ( .I(reorder_O2[22]), .ZN(n7365) );
  inv0d1 U9208 ( .I(reorder_O2[23]), .ZN(n7363) );
  inv0d1 U9209 ( .I(reorder_O2[25]), .ZN(n7355) );
  inv0d1 U9210 ( .I(reorder_O2[26]), .ZN(n7348) );
  inv0d1 U9211 ( .I(reorder_O2[28]), .ZN(n7325) );
  inv0d1 U9212 ( .I(reorder_O2[29]), .ZN(n7322) );
  inv0d1 U9213 ( .I(reorder_O2[31]), .ZN(n7307) );
  inv0d1 U9214 ( .I(reorder_O1[30]), .ZN(n7445) );
  inv0d1 U9215 ( .I(reorder_O1[0]), .ZN(n7558) );
  inv0d1 U9216 ( .I(reorder_O1[1]), .ZN(n7514) );
  inv0d1 U9217 ( .I(reorder_O1[2]), .ZN(n7448) );
  inv0d1 U9218 ( .I(reorder_O1[3]), .ZN(n7438) );
  inv0d1 U9219 ( .I(reorder_O1[4]), .ZN(n7432) );
  inv0d1 U9220 ( .I(reorder_O1[5]), .ZN(n7425) );
  inv0d1 U9221 ( .I(reorder_O1[6]), .ZN(n7424) );
  inv0d1 U9222 ( .I(reorder_O1[7]), .ZN(n7415) );
  inv0d1 U9223 ( .I(reorder_O1[8]), .ZN(n7414) );
  inv0d1 U9225 ( .I(reorder_O1[9]), .ZN(n7412) );
  inv0d1 U9226 ( .I(reorder_O1[10]), .ZN(n7553) );
  inv0d1 U9227 ( .I(reorder_O1[11]), .ZN(n7552) );
  inv0d1 U9228 ( .I(reorder_O1[12]), .ZN(n7549) );
  inv0d1 U9229 ( .I(reorder_O1[13]), .ZN(n7542) );
  inv0d1 U9230 ( .I(reorder_O1[14]), .ZN(n7538) );
  inv0d1 U9231 ( .I(reorder_O1[15]), .ZN(n7531) );
  inv0d1 U9232 ( .I(reorder_O1[16]), .ZN(n7525) );
  inv0d1 U9233 ( .I(reorder_O1[17]), .ZN(n7524) );
  inv0d1 U9234 ( .I(reorder_O1[18]), .ZN(n7520) );
  inv0d1 U9235 ( .I(reorder_O1[19]), .ZN(n7519) );
  inv0d1 U9236 ( .I(reorder_O1[20]), .ZN(n7510) );
  inv0d1 U9237 ( .I(reorder_O1[21]), .ZN(n7503) );
  inv0d1 U9238 ( .I(reorder_O1[22]), .ZN(n7497) );
  inv0d1 U9239 ( .I(reorder_O1[23]), .ZN(n7482) );
  inv0d1 U9240 ( .I(reorder_O1[24]), .ZN(n7476) );
  inv0d1 U9241 ( .I(reorder_O1[25]), .ZN(n7470) );
  inv0d1 U9242 ( .I(reorder_O1[26]), .ZN(n7467) );
  inv0d1 U9243 ( .I(reorder_O1[27]), .ZN(n7465) );
  inv0d1 U9244 ( .I(reorder_O1[28]), .ZN(n7451) );
  inv0d1 U9245 ( .I(reorder_O1[29]), .ZN(n7449) );
  inv0d1 U9246 ( .I(reorder_O1[31]), .ZN(n7441) );
  inv0d0 U9248 ( .I(N5027), .ZN(n2745) );
  inv0d0 U9249 ( .I(N5026), .ZN(n2746) );
  inv0d0 U9250 ( .I(N5028), .ZN(n2744) );
  inv0d0 U9251 ( .I(N5025), .ZN(n2747) );
  inv0d0 U9253 ( .I(N5024), .ZN(n2748) );
  nd02d1 U9254 ( .A1(n3597), .A2(n3598), .ZN(n12096) );
  nd02d1 U9255 ( .A1(n3599), .A2(n3600), .ZN(n12097) );
  nd02d1 U9256 ( .A1(n3601), .A2(n3602), .ZN(n12098) );
  nd02d1 U9257 ( .A1(n3603), .A2(n3604), .ZN(n12099) );
  nd02d1 U9259 ( .A1(n3605), .A2(n3606), .ZN(n12100) );
  nd02d1 U9260 ( .A1(n3611), .A2(n3612), .ZN(n12102) );
  nd02d1 U9261 ( .A1(n3613), .A2(n3614), .ZN(n12103) );
  nd02d1 U9262 ( .A1(n3615), .A2(n3616), .ZN(n12104) );
  inv0d0 U9263 ( .I(N5023), .ZN(n2749) );
  nd02d1 U9264 ( .A1(images_bus[2]), .A2(n477), .ZN(n417) );
  inv0d0 U9265 ( .I(n12130), .ZN(n6806) );
  inv0d0 U9266 ( .I(n12124), .ZN(n6901) );
  inv0d0 U9267 ( .I(N5022), .ZN(n2750) );
  nd02d1 U9268 ( .A1(n3628), .A2(n3629), .ZN(n12108) );
  nd02d1 U9269 ( .A1(n3630), .A2(n3631), .ZN(n12109) );
  nd02d1 U9270 ( .A1(n3632), .A2(n3633), .ZN(n12110) );
  nd02d1 U9271 ( .A1(n3634), .A2(n3635), .ZN(n12111) );
  nd02d1 U9272 ( .A1(n3636), .A2(n3637), .ZN(n12112) );
  nd02d1 U9273 ( .A1(n3638), .A2(n3639), .ZN(n12113) );
  nd02d1 U9274 ( .A1(n3644), .A2(n3645), .ZN(n12116) );
  nd02d1 U9275 ( .A1(n3640), .A2(n3641), .ZN(n12114) );
  nd02d1 U9277 ( .A1(n3642), .A2(n3643), .ZN(n12115) );
  inv0d0 U9278 ( .I(N5021), .ZN(n2751) );
  nd02d1 U9279 ( .A1(n2754), .A2(n3588), .ZN(n3579) );
  nd02d1 U9280 ( .A1(n3626), .A2(n3627), .ZN(n12107) );
  nd02d1 U9281 ( .A1(N3878), .A2(n949), .ZN(n3627) );
  nd02d1 U9282 ( .A1(n3624), .A2(n3625), .ZN(n12106) );
  nd02d1 U9283 ( .A1(N3877), .A2(n949), .ZN(n3625) );
  nd02d1 U9284 ( .A1(n3591), .A2(n3592), .ZN(n12094) );
  nd02d1 U9285 ( .A1(N3877), .A2(n949), .ZN(n3592) );
  nd02d1 U9286 ( .A1(n3595), .A2(n3596), .ZN(n12095) );
  nd02d1 U9287 ( .A1(N3878), .A2(n949), .ZN(n3596) );
  nd04d1 U9288 ( .A1(N5029), .A2(n4235), .A3(distance_ready), .A4(n4242), .ZN(
        n4240) );
  nd03d1 U9289 ( .A1(n493), .A2(n2774), .A3(hashes_ready), .ZN(n4237) );
  inv0d0 U9290 ( .I(N5020), .ZN(n2752) );
  nd03d1 U9292 ( .A1(distance_ready), .A2(N4760), .A3(hashes_ready), .ZN(n3676) );
  inv0d0 U9294 ( .I(n12169), .ZN(n4946) );
  inv0d0 U9295 ( .I(n12149), .ZN(n6466) );
  nd03d1 U9296 ( .A1(n2771), .A2(n4242), .A3(new_reference_is_done), .ZN(n4241) );
  an03d1 U9297 ( .A1(N5029), .A2(n4235), .A3(n4236), .Z(n4234) );
  inv0d0 U9298 ( .I(n12122), .ZN(n6922) );
  inv0d0 U9299 ( .I(n12132), .ZN(n6737) );
  inv0d0 U9300 ( .I(n12157), .ZN(n6235) );
  inv0d0 U9301 ( .I(n12168), .ZN(n4958) );
  inv0d0 U9302 ( .I(n12143), .ZN(n6547) );
  inv0d0 U9303 ( .I(n12120), .ZN(n6967) );
  nd02d1 U9304 ( .A1(N3187), .A2(n2772), .ZN(n3657) );
  inv0d0 U9305 ( .I(count_image[8]), .ZN(n2738) );
  inv0d0 U9306 ( .I(count_image[7]), .ZN(n2742) );
  inv0d0 U9307 ( .I(n12167), .ZN(n5354) );
  inv0d0 U9309 ( .I(n12128), .ZN(n6861) );
  inv0d0 U9310 ( .I(n12170), .ZN(n4698) );
  inv0d0 U9311 ( .I(n12148), .ZN(n6496) );
  inv0d0 U9312 ( .I(n12129), .ZN(n6818) );
  inv0d0 U9313 ( .I(n2726), .ZN(n2740) );
  inv0d0 U9314 ( .I(count_image[0]), .ZN(n2741) );
  inv0d0 U9316 ( .I(count_image[3]), .ZN(n2739) );
  inv0d0 U9317 ( .I(n12131), .ZN(n6795) );
  inv0d0 U9318 ( .I(n12165), .ZN(n5626) );
  inv0d0 U9319 ( .I(n12135), .ZN(n6664) );
  inv0d0 U9320 ( .I(n12140), .ZN(n6599) );
  inv0d0 U9321 ( .I(n12119), .ZN(n7062) );
  inv0d0 U9322 ( .I(n12151), .ZN(n6425) );
  inv0d0 U9325 ( .I(n12126), .ZN(n6890) );
  inv0d0 U9326 ( .I(n12146), .ZN(n6531) );
  inv0d0 U9327 ( .I(n12156), .ZN(n6279) );
  inv0d0 U9328 ( .I(n12127), .ZN(n6871) );
  inv0d0 U9329 ( .I(n12153), .ZN(n6383) );
  inv0d0 U9330 ( .I(n12172), .ZN(n4331) );
  inv0d0 U9331 ( .I(n12150), .ZN(n6437) );
  inv0d0 U9332 ( .I(n12133), .ZN(n6699) );
  inv0d0 U9333 ( .I(n12118), .ZN(n7153) );
  inv0d0 U9334 ( .I(n12138), .ZN(n6601) );
  inv0d0 U9335 ( .I(n12171), .ZN(n4416) );
  inv0d0 U9336 ( .I(n12161), .ZN(n6155) );
  inv0d0 U9337 ( .I(n12142), .ZN(n6556) );
  inv0d0 U9338 ( .I(n12136), .ZN(n6659) );
  inv0d0 U9339 ( .I(n12144), .ZN(n6544) );
  inv0d0 U9340 ( .I(n12164), .ZN(n5714) );
  inv0d0 U9341 ( .I(n12160), .ZN(n6157) );
  inv0d0 U9342 ( .I(n12147), .ZN(n6512) );
  inv0d0 U9343 ( .I(n12139), .ZN(n6600) );
  inv0d0 U9344 ( .I(n12125), .ZN(n6892) );
  inv0d0 U9345 ( .I(n12123), .ZN(n6908) );
  inv0d0 U9346 ( .I(n12159), .ZN(n6179) );
  inv0d0 U9347 ( .I(n12155), .ZN(n6324) );
  inv0d0 U9348 ( .I(n12154), .ZN(n6328) );
  inv0d0 U9349 ( .I(n12187), .ZN(\lt_82/A[5] ) );
  inv0d0 U9350 ( .I(n12141), .ZN(n6598) );
  inv0d0 U9351 ( .I(n12152), .ZN(n6423) );
  inv0d0 U9352 ( .I(n12134), .ZN(n6682) );
  inv0d0 U9353 ( .I(n12145), .ZN(n6543) );
  inv0d0 U9354 ( .I(n12166), .ZN(n5604) );
  inv0d0 U9355 ( .I(n12121), .ZN(n6931) );
  inv0d0 U9356 ( .I(n12173), .ZN(n4297) );
  inv0d0 U9357 ( .I(n12158), .ZN(n6212) );
  inv0d0 U9358 ( .I(n3661), .ZN(n2767) );
  inv0d0 U9360 ( .I(N29403), .ZN(n2780) );
  nr02d1 U9361 ( .A1(n2758), .A2(n12204), .ZN(n3794) );
  inv0d0 U9362 ( .I(images_bus[418]), .ZN(n6897) );
  inv0d0 U9363 ( .I(images_bus[434]), .ZN(n6732) );
  inv0d0 U9365 ( .I(n12137), .ZN(n6621) );
  inv0d0 U9366 ( .I(images_bus[484]), .ZN(n6596) );
  nr02d1 U9367 ( .A1(temp_new_reference[8]), .A2(n2758), .ZN(n4010) );
  inv0d0 U9368 ( .I(images_bus[32]), .ZN(n7260) );
  inv0d0 U9370 ( .I(images_bus[64]), .ZN(n7255) );
  inv0d0 U9371 ( .I(images_bus[210]), .ZN(n6776) );
  inv0d0 U9372 ( .I(images_bus[122]), .ZN(n6698) );
  inv0d0 U9373 ( .I(images_bus[132]), .ZN(n6638) );
  inv0d0 U9374 ( .I(images_bus[65]), .ZN(n5776) );
  inv0d0 U9377 ( .I(images_bus[19]), .ZN(n5113) );
  inv0d0 U9378 ( .I(images_bus[27]), .ZN(n4976) );
  inv0d0 U9379 ( .I(images_bus[133]), .ZN(n4727) );
  inv0d0 U9380 ( .I(n12162), .ZN(n6152) );
  inv0d0 U9381 ( .I(images_bus[94]), .ZN(n6199) );
  inv0d0 U9382 ( .I(images_bus[222]), .ZN(n6176) );
  inv0d0 U9383 ( .I(n12163), .ZN(n6147) );
  inv0d0 U9384 ( .I(images_bus[384]), .ZN(n7207) );
  inv0d0 U9385 ( .I(images_bus[282]), .ZN(n6676) );
  inv0d0 U9386 ( .I(images_bus[364]), .ZN(n6560) );
  inv0d0 U9387 ( .I(images_bus[404]), .ZN(n6523) );
  inv0d0 U9388 ( .I(images_bus[463]), .ZN(n5898) );
  inv0d0 U9389 ( .I(images_bus[380]), .ZN(n6443) );
  inv0d0 U9390 ( .I(n12188), .ZN(\lt_82/A[4] ) );
  inv0d0 U9391 ( .I(n4340), .ZN(n2763) );
  inv0d0 U9392 ( .I(n4336), .ZN(n2764) );
  inv0d0 U9393 ( .I(n4349), .ZN(n2761) );
  inv0d0 U9394 ( .I(n4332), .ZN(n2765) );
  inv0d0 U9395 ( .I(n4350), .ZN(n2760) );
  inv0d0 U9396 ( .I(n4344), .ZN(n2762) );
  inv0d0 U9397 ( .I(compare_in_progress), .ZN(n2787) );
  inv0d0 U9398 ( .I(n3669), .ZN(n2769) );
  inv0d0 U9399 ( .I(finish_flag), .ZN(n2772) );
  inv0d0 U9400 ( .I(n12174), .ZN(\add_0_root_add_1_root_add_98_3/A[3] ) );
  inv0d0 U9401 ( .I(hashes_ready), .ZN(n2776) );
  nd03d1 U9403 ( .A1(n2776), .A2(n2779), .A3(compare_in_progress), .ZN(n3685)
         );
  nd02d1 U9404 ( .A1(reading_compare), .A2(n2776), .ZN(n3656) );
  inv0d0 U9406 ( .I(reading_compare), .ZN(n2779) );
  inv0d0 U9407 ( .I(n12177), .ZN(\add_0_root_add_1_root_add_98_3/A[4] ) );
  inv0d0 U9408 ( .I(N3878), .ZN(n2789) );
  oai21d1 U9409 ( .B1(distance[8]), .B2(n12091), .A(n1418), .ZN(N5029) );
  nd04d1 U9410 ( .A1(n2784), .A2(n2739), .A3(n4377), .A4(n4378), .ZN(N26489)
         );
  inv0d0 U9412 ( .I(n1407), .ZN(n1419) );
  inv0d0 U9413 ( .I(count_image[2]), .ZN(n2784) );
  inv0d0 U9414 ( .I(n12178), .ZN(\add_0_root_add_1_root_add_98_3/A[5] ) );
  inv0d0 U9415 ( .I(n12179), .ZN(\add_0_root_add_1_root_add_98_3/A[6] ) );
  inv0d0 U9416 ( .I(N3877), .ZN(n2788) );
  inv0d0 U9417 ( .I(n12180), .ZN(\add_0_root_add_1_root_add_98_3/A[7] ) );
  nd02d1 U9418 ( .A1(reading_current), .A2(n2776), .ZN(n3654) );
  inv0d0 U9421 ( .I(n12181), .ZN(\add_0_root_add_1_root_add_98_3/A[8] ) );
  inv0d0 U9423 ( .I(n12182), .ZN(\add_0_root_add_1_root_add_98_3/A[9] ) );
  nr02d1 U9424 ( .A1(n12208), .A2(N3234), .ZN(n4212) );
  nr02d1 U9425 ( .A1(N3234), .A2(N3235), .ZN(n4192) );
  nr02d1 U9426 ( .A1(n12209), .A2(N3235), .ZN(n4221) );
  nr02d1 U9427 ( .A1(temp_new_reference[5]), .A2(n12205), .ZN(n3796) );
  nr02d1 U9428 ( .A1(temp_new_reference[7]), .A2(temp_new_reference[6]), .ZN(
        n3948) );
  nr02d1 U9429 ( .A1(temp_new_reference[7]), .A2(n12206), .ZN(n3884) );
  nr02d1 U9430 ( .A1(n12209), .A2(n12208), .ZN(n4197) );
  nr02d1 U9431 ( .A1(n12205), .A2(n12207), .ZN(n3825) );
  inv0d0 U9433 ( .I(n12183), .ZN(\add_0_root_add_1_root_add_98_3/A[10] ) );
  inv0d0 U9437 ( .I(distance_ready), .ZN(n2778) );
  inv0d0 U9438 ( .I(n12207), .ZN(n2785) );
  inv0d0 U9441 ( .I(n12206), .ZN(n2786) );
  inv0d0 U9442 ( .I(n12184), .ZN(\add_0_root_add_1_root_add_98_3/A[11] ) );
  nr02d1 U9443 ( .A1(n3697), .A2(n3698), .ZN(n3696) );
  inv0d0 U9444 ( .I(new_reference_is_done), .ZN(n2782) );
  inv0d0 U9445 ( .I(images_bus[399]), .ZN(n5906) );
  inv0d0 U9446 ( .I(images_bus[195]), .ZN(n5276) );
  inv0d0 U9448 ( .I(images_bus[271]), .ZN(n5933) );
  inv0d0 U9450 ( .I(images_bus[204]), .ZN(n6571) );
  inv0d0 U9451 ( .I(images_bus[444]), .ZN(n6428) );
  inv0d0 U9453 ( .I(images_bus[13]), .ZN(n4608) );
  inv0d0 U9454 ( .I(images_bus[407]), .ZN(n5806) );
  inv0d0 U9455 ( .I(images_bus[119]), .ZN(n5855) );
  inv0d0 U9456 ( .I(images_bus[207]), .ZN(n5944) );
  inv0d0 U9457 ( .I(images_bus[319]), .ZN(n6098) );
  inv0d0 U9458 ( .I(images_bus[416]), .ZN(n7205) );
  inv0d0 U9459 ( .I(images_bus[303]), .ZN(n5931) );
  inv0d0 U9460 ( .I(images_bus[264]), .ZN(n7152) );
  inv0d0 U9461 ( .I(images_bus[363]), .ZN(n5146) );
  inv0d0 U9462 ( .I(images_bus[325]), .ZN(n4663) );
  inv0d0 U9463 ( .I(images_bus[104]), .ZN(n7176) );
  inv0d0 U9464 ( .I(images_bus[203]), .ZN(n5186) );
  inv0d0 U9465 ( .I(images_bus[139]), .ZN(n5194) );
  inv0d0 U9466 ( .I(images_bus[414]), .ZN(n6160) );
  inv0d0 U9467 ( .I(images_bus[343]), .ZN(n5825) );
  inv0d0 U9468 ( .I(images_bus[79]), .ZN(n5958) );
  inv0d0 U9469 ( .I(images_bus[339]), .ZN(n5046) );
  inv0d0 U9470 ( .I(images_bus[223]), .ZN(n6115) );
  inv0d0 U9471 ( .I(images_bus[403]), .ZN(n5034) );
  inv0d0 U9472 ( .I(images_bus[408]), .ZN(n6993) );
  inv0d0 U9473 ( .I(images_bus[423]), .ZN(n5980) );
  inv0d0 U9474 ( .I(images_bus[163]), .ZN(n5278) );
  inv0d0 U9475 ( .I(images_bus[359]), .ZN(n5988) );
  inv0d0 U9476 ( .I(images_bus[152]), .ZN(n7023) );
  inv0d0 U9477 ( .I(images_bus[496]), .ZN(n7050) );
  inv0d0 U9478 ( .I(images_bus[141]), .ZN(n4491) );
  inv0d0 U9479 ( .I(images_bus[55]), .ZN(n5862) );
  inv0d0 U9481 ( .I(images_bus[415]), .ZN(n6084) );
  inv0d0 U9482 ( .I(images_bus[297]), .ZN(n5636) );
  inv0d0 U9483 ( .I(images_bus[495]), .ZN(n5894) );
  inv0d0 U9484 ( .I(images_bus[253]), .ZN(n3577) );
  inv0d0 U9485 ( .I(images_bus[453]), .ZN(n4635) );
  inv0d0 U9486 ( .I(images_bus[96]), .ZN(n7251) );
  inv0d0 U9487 ( .I(images_bus[103]), .ZN(n6056) );
  inv0d0 U9489 ( .I(images_bus[176]), .ZN(n7081) );
  inv0d0 U9491 ( .I(images_bus[140]), .ZN(n6575) );
  inv0d0 U9492 ( .I(images_bus[105]), .ZN(n5689) );
  inv0d0 U9493 ( .I(images_bus[211]), .ZN(n5068) );
  inv0d0 U9494 ( .I(images_bus[405]), .ZN(n4302) );
  inv0d0 U9495 ( .I(images_bus[168]), .ZN(n7166) );
  inv0d0 U9496 ( .I(images_bus[323]), .ZN(n5254) );
  inv0d0 U9497 ( .I(images_bus[235]), .ZN(n5173) );
  inv0d0 U9498 ( .I(images_bus[182]), .ZN(n6259) );
  inv0d0 U9500 ( .I(images_bus[39]), .ZN(n6070) );
  inv0d0 U9501 ( .I(images_bus[287]), .ZN(n6100) );
  inv0d0 U9502 ( .I(images_bus[208]), .ZN(n7079) );
  inv0d0 U9505 ( .I(images_bus[324]), .ZN(n6606) );
  inv0d0 U9507 ( .I(images_bus[279]), .ZN(n5834) );
  inv0d0 U9508 ( .I(images_bus[345]), .ZN(n5397) );
  inv0d0 U9509 ( .I(images_bus[111]), .ZN(n5957) );
  inv0d0 U9510 ( .I(images_bus[67]), .ZN(n5298) );
  inv0d0 U9512 ( .I(images_bus[101]), .ZN(n4745) );
  inv0d0 U9513 ( .I(images_bus[352]), .ZN(n7222) );
  inv0d0 U9515 ( .I(images_bus[413]), .ZN(n3129) );
  inv0d0 U9516 ( .I(images_bus[483]), .ZN(n5221) );
  inv0d0 U9517 ( .I(images_bus[437]), .ZN(n4300) );
  inv0d0 U9518 ( .I(images_bus[500]), .ZN(n6508) );
  inv0d0 U9519 ( .I(images_bus[44]), .ZN(n6589) );
  inv0d0 U9520 ( .I(images_bus[41]), .ZN(n5704) );
  inv0d0 U9522 ( .I(images_bus[131]), .ZN(n5281) );
  inv0d0 U9523 ( .I(images_bus[75]), .ZN(n5204) );
  inv0d0 U9524 ( .I(images_bus[88]), .ZN(n7042) );
  inv0d0 U9527 ( .I(images_bus[293]), .ZN(n4675) );
  inv0d0 U9528 ( .I(images_bus[455]), .ZN(n5979) );
  inv0d0 U9529 ( .I(images_bus[221]), .ZN(n3619) );
  inv0d0 U9530 ( .I(images_bus[224]), .ZN(n7242) );
  inv0d0 U9531 ( .I(images_bus[112]), .ZN(n7097) );
  inv0d0 U9532 ( .I(images_bus[328]), .ZN(n7136) );
  inv0d0 U9533 ( .I(images_bus[199]), .ZN(n6038) );
  inv0d0 U9535 ( .I(images_bus[429]), .ZN(n4406) );
  inv0d0 U9536 ( .I(images_bus[169]), .ZN(n5676) );
  inv0d0 U9537 ( .I(images_bus[134]), .ZN(n6397) );
  inv0d0 U9539 ( .I(images_bus[307]), .ZN(n5049) );
  inv0d0 U9540 ( .I(images_bus[31]), .ZN(n6146) );
  inv0d0 U9542 ( .I(images_bus[61]), .ZN(n4222) );
  inv0d0 U9543 ( .I(images_bus[69]), .ZN(n4751) );
  inv0d0 U9544 ( .I(images_bus[504]), .ZN(n6979) );
  inv0d0 U9545 ( .I(images_bus[391]), .ZN(n5982) );
  inv0d0 U9546 ( .I(images_bus[198]), .ZN(n6390) );
  inv0d0 U9548 ( .I(images_bus[229]), .ZN(n4691) );
  inv0d0 U9550 ( .I(images_bus[175]), .ZN(n5949) );
  inv0d0 U9551 ( .I(images_bus[243]), .ZN(n5063) );
  inv0d0 U9552 ( .I(images_bus[471]), .ZN(n5798) );
  inv0d0 U9553 ( .I(images_bus[299]), .ZN(n5164) );
  inv0d0 U9554 ( .I(images_bus[68]), .ZN(n6641) );
  inv0d0 U9555 ( .I(images_bus[120]), .ZN(n7034) );
  inv0d0 U9556 ( .I(images_bus[304]), .ZN(n7072) );
  inv0d0 U9557 ( .I(images_bus[37]), .ZN(n4754) );
  inv0d0 U9558 ( .I(images_bus[424]), .ZN(n7121) );
  inv0d0 U9559 ( .I(images_bus[144]), .ZN(n7093) );
  inv0d0 U9560 ( .I(images_bus[42]), .ZN(n6884) );
  inv0d0 U9561 ( .I(images_bus[196]), .ZN(n6628) );
  inv0d0 U9562 ( .I(images_bus[381]), .ZN(n3138) );
  inv0d0 U9563 ( .I(images_bus[107]), .ZN(n5203) );
  inv0d0 U9565 ( .I(images_bus[340]), .ZN(n6529) );
  inv0d0 U9566 ( .I(images_bus[443]), .ZN(n4894) );
  inv0d0 U9567 ( .I(images_bus[315]), .ZN(n4939) );
  inv0d0 U9568 ( .I(images_bus[288]), .ZN(n7237) );
  inv0d0 U9569 ( .I(images_bus[73]), .ZN(n5691) );
  inv0d0 U9570 ( .I(images_bus[367]), .ZN(n5920) );
  inv0d0 U9571 ( .I(images_bus[486]), .ZN(n6356) );
  inv0d0 U9573 ( .I(images_bus[255]), .ZN(n6113) );
  inv0d0 U9574 ( .I(images_bus[346]), .ZN(n6670) );
  inv0d0 U9576 ( .I(images_bus[173]), .ZN(n4464) );
  inv0d0 U9578 ( .I(images_bus[427]), .ZN(n5136) );
  inv0d0 U9579 ( .I(images_bus[375]), .ZN(n5818) );
  inv0d0 U9580 ( .I(images_bus[344]), .ZN(n6998) );
  inv0d0 U9581 ( .I(images_bus[440]), .ZN(n6990) );
  inv0d0 U9582 ( .I(images_bus[333]), .ZN(n4427) );
  inv0d0 U9583 ( .I(images_bus[177]), .ZN(n5558) );
  inv0d0 U9584 ( .I(images_bus[417]), .ZN(n5728) );
  inv0d0 U9588 ( .I(images_bus[167]), .ZN(n6039) );
  inv0d0 U9589 ( .I(images_bus[289]), .ZN(n5738) );
  inv0d0 U9590 ( .I(images_bus[379]), .ZN(n4902) );
  inv0d0 U9591 ( .I(images_bus[231]), .ZN(n6025) );
  inv0d0 U9593 ( .I(images_bus[183]), .ZN(n5846) );
  inv0d0 U9594 ( .I(images_bus[143]), .ZN(n5952) );
  inv0d0 U9596 ( .I(images_bus[274]), .ZN(n6753) );
  inv0d0 U9597 ( .I(images_bus[80]), .ZN(n7104) );
  inv0d0 U9598 ( .I(images_bus[311]), .ZN(n5826) );
  inv0d0 U9599 ( .I(images_bus[436]), .ZN(n6519) );
  inv0d0 U9601 ( .I(images_bus[85]), .ZN(n4326) );
  inv0d0 U9602 ( .I(images_bus[438]), .ZN(n6218) );
  inv0d0 U9603 ( .I(images_bus[357]), .ZN(n4653) );
  inv0d0 U9604 ( .I(images_bus[419]), .ZN(n5235) );
  inv0d0 U9605 ( .I(images_bus[251]), .ZN(n4948) );
  inv0d0 U9606 ( .I(images_bus[159]), .ZN(n6123) );
  inv0d0 U9607 ( .I(images_bus[292]), .ZN(n6613) );
  inv0d0 U9608 ( .I(images_bus[239]), .ZN(n5937) );
  inv0d0 U9610 ( .I(images_bus[347]), .ZN(n4915) );
  inv0d0 U9612 ( .I(images_bus[127]), .ZN(n6133) );
  inv0d0 U9613 ( .I(images_bus[87]), .ZN(n5858) );
  inv0d0 U9614 ( .I(images_bus[247]), .ZN(n5835) );
  inv0d0 U9615 ( .I(images_bus[145]), .ZN(n5573) );
  inv0d0 U9616 ( .I(images_bus[326]), .ZN(n6371) );
  inv0d0 U9617 ( .I(images_bus[327]), .ZN(n6004) );
  inv0d0 U9618 ( .I(images_bus[448]), .ZN(n7194) );
  inv0d0 U9619 ( .I(images_bus[76]), .ZN(n6586) );
  inv0d0 U9620 ( .I(images_bus[188]), .ZN(n6481) );
  inv0d0 U9621 ( .I(images_bus[313]), .ZN(n5405) );
  inv0d0 U9622 ( .I(images_bus[268]), .ZN(n6566) );
  inv0d0 U9623 ( .I(images_bus[220]), .ZN(n6475) );
  inv0d0 U9625 ( .I(images_bus[209]), .ZN(n5548) );
  inv0d0 U9629 ( .I(images_bus[435]), .ZN(n5003) );
  inv0d0 U9630 ( .I(images_bus[425]), .ZN(n5617) );
  inv0d0 U9631 ( .I(images_bus[295]), .ZN(n6007) );
  inv0d0 U9632 ( .I(images_bus[262]), .ZN(n6388) );
  inv0d0 U9633 ( .I(images_bus[51]), .ZN(n5110) );
  inv0d0 U9634 ( .I(images_bus[123]), .ZN(n4965) );
  inv0d0 U9635 ( .I(images_bus[406]), .ZN(n6225) );
  inv0d0 U9636 ( .I(images_bus[237]), .ZN(n4451) );
  inv0d0 U9637 ( .I(images_bus[136]), .ZN(n7173) );
  inv0d0 U9638 ( .I(images_bus[396]), .ZN(n6558) );
  inv0d0 U9639 ( .I(images_bus[309]), .ZN(n4307) );
  inv0d0 U9640 ( .I(images_bus[275]), .ZN(n5060) );
  inv0d0 U9641 ( .I(images_bus[296]), .ZN(n7150) );
  inv0d0 U9642 ( .I(images_bus[464]), .ZN(n7057) );
  inv0d0 U9643 ( .I(images_bus[371]), .ZN(n5043) );
  inv0d0 U9644 ( .I(images_bus[15]), .ZN(n5964) );
  inv0d0 U9646 ( .I(images_bus[479]), .ZN(n6074) );
  inv0d0 U9647 ( .I(images_bus[45]), .ZN(n4512) );
  inv0d0 U9648 ( .I(images_bus[459]), .ZN(n5126) );
  inv0d0 U9649 ( .I(images_bus[205]), .ZN(n4459) );
  inv0d0 U9650 ( .I(images_bus[216]), .ZN(n7019) );
  inv0d0 U9652 ( .I(images_bus[329]), .ZN(n5633) );
  inv0d0 U9653 ( .I(images_bus[97]), .ZN(n5775) );
  inv0d0 U9654 ( .I(images_bus[89]), .ZN(n5456) );
  inv0d0 U9656 ( .I(images_bus[121]), .ZN(n5447) );
  inv0d0 U9657 ( .I(images_bus[108]), .ZN(n6576) );
  inv0d0 U9658 ( .I(images_bus[421]), .ZN(n4640) );
  inv0d0 U9660 ( .I(images_bus[451]), .ZN(n5231) );
  inv0d0 U9661 ( .I(images_bus[387]), .ZN(n5242) );
  inv0d0 U9662 ( .I(images_bus[373]), .ZN(n4304) );
  inv0d0 U9663 ( .I(images_bus[472]), .ZN(n6982) );
  inv0d0 U9664 ( .I(images_bus[130]), .ZN(n6946) );
  inv0d0 U9665 ( .I(images_bus[505]), .ZN(n5320) );
  inv0d0 U9666 ( .I(images_bus[149]), .ZN(n4319) );
  inv0d0 U9667 ( .I(images_bus[125]), .ZN(n3986) );
  inv0d0 U9668 ( .I(images_bus[109]), .ZN(n4493) );
  inv0d0 U9669 ( .I(images_bus[259]), .ZN(n5266) );
  inv0d0 U9670 ( .I(images_bus[457]), .ZN(n5607) );
  inv0d0 U9671 ( .I(images_bus[477]), .ZN(n2819) );
  inv0d0 U9675 ( .I(images_bus[369]), .ZN(n5523) );
  inv0d0 U9676 ( .I(images_bus[280]), .ZN(n7016) );
  inv0d0 U9677 ( .I(images_bus[213]), .ZN(n4314) );
  inv0d0 U9678 ( .I(images_bus[503]), .ZN(n5797) );
  inv0d0 U9679 ( .I(images_bus[74]), .ZN(n6882) );
  inv0d0 U9680 ( .I(images_bus[219]), .ZN(n4951) );
  inv0d0 U9682 ( .I(images_bus[317]), .ZN(n3331) );
  inv0d0 U9683 ( .I(images_bus[411]), .ZN(n4900) );
  inv0d0 U9684 ( .I(images_bus[382]), .ZN(n6162) );
  inv0d0 U9685 ( .I(images_bus[161]), .ZN(n5762) );
  inv0d0 U9686 ( .I(images_bus[291]), .ZN(n5265) );
  inv0d0 U9688 ( .I(images_bus[474]), .ZN(n6655) );
  inv0d0 U9689 ( .I(images_bus[305]), .ZN(n5531) );
  inv0d0 U9690 ( .I(images_bus[240]), .ZN(n7076) );
  inv0d0 U9691 ( .I(images_bus[321]), .ZN(n5737) );
  inv0d0 U9692 ( .I(images_bus[1]), .ZN(n5785) );
  inv0d0 U9693 ( .I(images_bus[81]), .ZN(n5581) );
  inv0d0 U9694 ( .I(images_bus[227]), .ZN(n5268) );
  inv0d0 U9695 ( .I(images_bus[25]), .ZN(n5466) );
  inv0d0 U9696 ( .I(images_bus[84]), .ZN(n6548) );
  inv0d0 U9698 ( .I(images_bus[58]), .ZN(n6701) );
  inv0d0 U9699 ( .I(images_bus[439]), .ZN(n5802) );
  inv0d0 U9700 ( .I(images_bus[215]), .ZN(n5839) );
  inv0d0 U9701 ( .I(images_bus[35]), .ZN(n5312) );
  inv0d0 U9702 ( .I(images_bus[312]), .ZN(n7006) );
  inv0d0 U9703 ( .I(images_bus[91]), .ZN(n4973) );
  inv0d0 U9708 ( .I(images_bus[497]), .ZN(n5470) );
  inv0d0 U9709 ( .I(images_bus[241]), .ZN(n5542) );
  inv0d0 U9710 ( .I(images_bus[447]), .ZN(n6083) );
  inv0d0 U9711 ( .I(images_bus[286]), .ZN(n6173) );
  inv0d0 U9712 ( .I(images_bus[449]), .ZN(n5727) );
  inv0d0 U9714 ( .I(images_bus[157]), .ZN(n3903) );
  inv0d0 U9715 ( .I(images_bus[395]), .ZN(n5145) );
  inv0d0 U9717 ( .I(images_bus[254]), .ZN(n6174) );
  inv0d0 U9718 ( .I(images_bus[214]), .ZN(n6250) );
  inv0d0 U9719 ( .I(images_bus[14]), .ZN(n6355) );
  inv0d0 U9720 ( .I(images_bus[450]), .ZN(n6894) );
  inv0d0 U9721 ( .I(images_bus[488]), .ZN(n7115) );
  inv0d0 U9722 ( .I(images_bus[277]), .ZN(n4311) );
  inv0d0 U9724 ( .I(images_bus[389]), .ZN(n4649) );
  inv0d0 U9725 ( .I(images_bus[469]), .ZN(n4298) );
  inv0d0 U9732 ( .I(images_bus[390]), .ZN(n6366) );
  inv0d0 U9733 ( .I(images_bus[57]), .ZN(n5459) );
  inv0d0 U9734 ( .I(images_bus[162]), .ZN(n6938) );
  inv0d0 U9735 ( .I(images_bus[300]), .ZN(n6565) );
  inv0d0 U9736 ( .I(images_bus[487]), .ZN(n5968) );
  inv0d0 U9738 ( .I(images_bus[24]), .ZN(n7047) );
  inv0d0 U9739 ( .I(images_bus[160]), .ZN(n7244) );
  inv0d0 U9740 ( .I(images_bus[171]), .ZN(n5189) );
  inv0d0 U9741 ( .I(images_bus[454]), .ZN(n6358) );
  inv0d0 U9742 ( .I(images_bus[355]), .ZN(n5249) );
  inv0d0 U9743 ( .I(images_bus[281]), .ZN(n5410) );
  inv0d0 U9744 ( .I(images_bus[86]), .ZN(n6268) );
  inv0d0 U9746 ( .I(images_bus[181]), .ZN(n4316) );
  inv0d0 U9747 ( .I(images_bus[358]), .ZN(n6368) );
  inv0d0 U9748 ( .I(images_bus[322]), .ZN(n6919) );
  inv0d0 U9749 ( .I(images_bus[402]), .ZN(n6736) );
  inv0d0 U9750 ( .I(images_bus[494]), .ZN(n6276) );
  inv0d0 U9751 ( .I(images_bus[147]), .ZN(n5098) );
  inv0d0 U9752 ( .I(images_bus[99]), .ZN(n5284) );
  inv0d0 U9753 ( .I(images_bus[166]), .ZN(n6395) );
  inv0d0 U9755 ( .I(images_bus[492]), .ZN(n6553) );
  inv0d0 U9756 ( .I(images_bus[93]), .ZN(n4119) );
  inv0d0 U9757 ( .I(images_bus[17]), .ZN(n5591) );
  inv0d0 U9758 ( .I(images_bus[341]), .ZN(n4306) );
  inv0d0 U9759 ( .I(images_bus[298]), .ZN(n6842) );
  inv0d0 U9760 ( .I(images_bus[431]), .ZN(n5902) );
  inv0d0 U9761 ( .I(images_bus[267]), .ZN(n5168) );
  inv0d0 U9762 ( .I(images_bus[400]), .ZN(n7066) );
  inv0d0 U9765 ( .I(images_bus[409]), .ZN(n5355) );
  inv0d0 U9766 ( .I(images_bus[460]), .ZN(n6555) );
  inv0d0 U9768 ( .I(images_bus[11]), .ZN(n5220) );
  inv0d0 U9769 ( .I(images_bus[155]), .ZN(n4959) );
  inv0d0 U9771 ( .I(images_bus[401]), .ZN(n5506) );
  inv0d0 U9772 ( .I(images_bus[465]), .ZN(n5484) );
  inv0d0 U9773 ( .I(images_bus[192]), .ZN(n7243) );
  inv0d0 U9774 ( .I(images_bus[48]), .ZN(n7105) );
  inv0d0 U9775 ( .I(images_bus[21]), .ZN(n4342) );
  inv0d0 U9778 ( .I(images_bus[164]), .ZN(n6630) );
  inv0d0 U9779 ( .I(images_bus[137]), .ZN(n5684) );
  inv0d0 U9781 ( .I(images_bus[485]), .ZN(n4633) );
  inv0d0 U9782 ( .I(images_bus[376]), .ZN(n6997) );
  inv0d0 U9784 ( .I(images_bus[7]), .ZN(n6072) );
  inv0d0 U9786 ( .I(images_bus[28]), .ZN(n6507) );
  inv0d0 U9787 ( .I(images_bus[77]), .ZN(n4503) );
  inv0d0 U9788 ( .I(images_bus[29]), .ZN(n4292) );
  inv0d0 U9789 ( .I(images_bus[2]), .ZN(n6975) );
  inv0d0 U9790 ( .I(images_bus[338]), .ZN(n6747) );
  inv0d0 U9791 ( .I(images_bus[233]), .ZN(n5648) );
  inv0d0 U9792 ( .I(images_bus[129]), .ZN(n5768) );
  inv0d0 U9793 ( .I(images_bus[249]), .ZN(n5426) );
  inv0d0 U9794 ( .I(images_bus[353]), .ZN(n5732) );
  inv0d0 U9795 ( .I(images_bus[115]), .ZN(n5104) );
  inv0d0 U9796 ( .I(images_bus[201]), .ZN(n5669) );
  inv0d0 U9797 ( .I(images_bus[200]), .ZN(n7155) );
  inv0d0 U9798 ( .I(images_bus[165]), .ZN(n4703) );
  inv0d0 U9799 ( .I(images_bus[475]), .ZN(n4890) );
  inv0d0 U9800 ( .I(images_bus[276]), .ZN(n6533) );
  inv0d0 U9801 ( .I(images_bus[135]), .ZN(n6051) );
  inv0d0 U9802 ( .I(images_bus[335]), .ZN(n5927) );
  inv0d0 U9803 ( .I(images_bus[445]), .ZN(n2915) );
  inv0d0 U9804 ( .I(images_bus[433]), .ZN(n5494) );
  inv0d0 U9805 ( .I(images_bus[331]), .ZN(n5156) );
  inv0d0 U9807 ( .I(images_bus[70]), .ZN(n6403) );
  inv0d0 U9809 ( .I(images_bus[40]), .ZN(n7183) );
  inv0d0 U9810 ( .I(images_bus[71]), .ZN(n6061) );
  inv0d0 U9811 ( .I(images_bus[490]), .ZN(n6817) );
  inv0d0 U9812 ( .I(images_bus[225]), .ZN(n5747) );
  inv0d0 U9813 ( .I(images_bus[20]), .ZN(n6552) );
  inv0d0 U9814 ( .I(images_bus[336]), .ZN(n7069) );
  inv0d0 U9815 ( .I(images_bus[368]), .ZN(n7067) );
  inv0d0 U9818 ( .I(images_bus[82]), .ZN(n6805) );
  inv0d0 U9819 ( .I(images_bus[473]), .ZN(n5322) );
  inv0d0 U9821 ( .I(images_bus[153]), .ZN(n5440) );
  inv0d0 U9822 ( .I(images_bus[269]), .ZN(n4450) );
  inv0d0 U9823 ( .I(images_bus[189]), .ZN(n3814) );
  inv0d0 U9824 ( .I(images_bus[194]), .ZN(n6934) );
  inv0d0 U9825 ( .I(images_bus[278]), .ZN(n6242) );
  inv0d0 U9826 ( .I(images_bus[59]), .ZN(n4974) );
  inv0d0 U9827 ( .I(images_bus[245]), .ZN(n4313) );
  inv0d0 U9828 ( .I(images_bus[493]), .ZN(n4393) );
  inv0d0 U9829 ( .I(images_bus[72]), .ZN(n7182) );
  inv0d0 U9830 ( .I(images_bus[461]), .ZN(n4397) );
  inv0d0 U9831 ( .I(images_bus[184]), .ZN(n7022) );
  inv0d0 U9832 ( .I(images_bus[481]), .ZN(n5715) );
  inv0d0 U9833 ( .I(images_bus[467]), .ZN(n4984) );
  inv0d0 U9834 ( .I(images_bus[285]), .ZN(n3478) );
  inv0d0 U9835 ( .I(images_bus[113]), .ZN(n5575) );
  inv0d0 U9836 ( .I(images_bus[128]), .ZN(n7245) );
  inv0d0 U9837 ( .I(images_bus[158]), .ZN(n6185) );
  inv0d0 U9839 ( .I(images_bus[244]), .ZN(n6538) );
  inv0d0 U9840 ( .I(images_bus[351]), .ZN(n6097) );
  inv0d0 U9842 ( .I(images_bus[22]), .ZN(n6273) );
  inv0d0 U9843 ( .I(images_bus[185]), .ZN(n5434) );
  inv0d0 U9844 ( .I(images_bus[334]), .ZN(n6297) );
  inv0d0 U9845 ( .I(images_bus[393]), .ZN(n5625) );
  inv0d0 U9850 ( .I(images_bus[316]), .ZN(n6455) );
  inv0d0 U9851 ( .I(images_bus[332]), .ZN(n6562) );
  inv0d0 U9852 ( .I(images_bus[350]), .ZN(n6166) );
  inv0d0 U9853 ( .I(images_bus[456]), .ZN(n7117) );
  inv0d0 U9854 ( .I(images_bus[320]), .ZN(n7232) );
  inv0d0 U9855 ( .I(images_bus[47]), .ZN(n5959) );
  inv0d0 U9857 ( .I(images_bus[248]), .ZN(n7017) );
  inv0d0 U9859 ( .I(images_bus[349]), .ZN(n3268) );
  inv0d0 U9860 ( .I(images_bus[117]), .ZN(n4321) );
  inv0d0 U9861 ( .I(images_bus[301]), .ZN(n4436) );
  inv0d0 U9862 ( .I(images_bus[272]), .ZN(n7075) );
  inv0d0 U9863 ( .I(images_bus[398]), .ZN(n6291) );
  inv0d0 U9864 ( .I(images_bus[236]), .ZN(n6567) );
  inv0d0 U9865 ( .I(images_bus[257]), .ZN(n5746) );
  inv0d0 U9866 ( .I(images_bus[179]), .ZN(n5079) );
  inv0d0 U9867 ( .I(images_bus[98]), .ZN(n6948) );
  inv0d0 U9868 ( .I(images_bus[56]), .ZN(n7045) );
  inv0d0 U9869 ( .I(images_bus[43]), .ZN(n5205) );
  inv0d0 U9870 ( .I(images_bus[430]), .ZN(n6287) );
  inv0d0 U9871 ( .I(images_bus[126]), .ZN(n6189) );
  inv0d0 U9873 ( .I(images_bus[365]), .ZN(n4419) );
  inv0d0 U9874 ( .I(images_bus[83]), .ZN(n5106) );
  inv0d0 U9876 ( .I(images_bus[49]), .ZN(n5585) );
  inv0d0 U9877 ( .I(images_bus[102]), .ZN(n6400) );
  inv0d0 U9878 ( .I(images_bus[366]), .ZN(n6293) );
  inv0d0 U9879 ( .I(images_bus[491]), .ZN(n5118) );
  inv0d0 U9880 ( .I(images_bus[38]), .ZN(n6411) );
  inv0d0 U9882 ( .I(images_bus[374]), .ZN(n6229) );
  inv0d0 U9883 ( .I(images_bus[191]), .ZN(n6119) );
  inv0d0 U9884 ( .I(images_bus[154]), .ZN(n6693) );
  inv0d0 U9885 ( .I(images_bus[310]), .ZN(n6240) );
  inv0d0 U9886 ( .I(images_bus[193]), .ZN(n5749) );
  inv0d0 U9887 ( .I(images_bus[499]), .ZN(n4980) );
  inv0d0 U9889 ( .I(images_bus[6]), .ZN(n6413) );
  inv0d0 U9891 ( .I(images_bus[242]), .ZN(n6759) );
  inv0d0 U9892 ( .I(images_bus[230]), .ZN(n6389) );
  inv0d0 U9893 ( .I(images_bus[156]), .ZN(n6484) );
  inv0d0 U9894 ( .I(images_bus[442]), .ZN(n6658) );
  inv0d0 U9895 ( .I(images_bus[256]), .ZN(n7240) );
  inv0d0 U9896 ( .I(images_bus[170]), .ZN(n6866) );
  inv0d0 U9897 ( .I(images_bus[507]), .ZN(n4886) );
  inv0d0 U9898 ( .I(images_bus[217]), .ZN(n5431) );
  inv0d0 U9899 ( .I(images_bus[265]), .ZN(n5644) );
  inv0d0 U9900 ( .I(images_bus[377]), .ZN(n5370) );
  inv0d0 U9901 ( .I(images_bus[480]), .ZN(n7188) );
  inv0d0 U9902 ( .I(images_bus[502]), .ZN(n6209) );
  inv0d0 U9903 ( .I(images_bus[16]), .ZN(n7109) );
  inv0d0 U9904 ( .I(images_bus[36]), .ZN(n6646) );
  inv0d0 U9905 ( .I(images_bus[314]), .ZN(n6675) );
  inv0d0 U9906 ( .I(images_bus[337]), .ZN(n5527) );
  inv0d0 U9907 ( .I(images_bus[151]), .ZN(n5851) );
  inv0d0 U9908 ( .I(images_bus[142]), .ZN(n6330) );
  inv0d0 U9909 ( .I(images_bus[63]), .ZN(n6140) );
  inv0d0 U9910 ( .I(images_bus[4]), .ZN(n6653) );
  inv0d0 U9911 ( .I(images_bus[385]), .ZN(n5730) );
  inv0d0 U9913 ( .I(images_bus[258]), .ZN(n6923) );
  inv0d0 U9914 ( .I(images_bus[263]), .ZN(n6024) );
  inv0d0 U9915 ( .I(images_bus[252]), .ZN(n6469) );
  inv0d0 U9919 ( .I(images_bus[18]), .ZN(n6813) );
  inv0d0 U9921 ( .I(images_bus[12]), .ZN(n6590) );
  inv0d0 U9922 ( .I(images_bus[234]), .ZN(n6855) );
  inv0d0 U9923 ( .I(images_bus[266]), .ZN(n6849) );
  inv0d0 U9924 ( .I(images_bus[150]), .ZN(n6264) );
  inv0d0 U9925 ( .I(images_bus[270]), .ZN(n6305) );
  inv0d0 U9926 ( .I(images_bus[260]), .ZN(n6618) );
  inv0d0 U9927 ( .I(images_bus[178]), .ZN(n6777) );
  inv0d0 U9928 ( .I(images_bus[106]), .ZN(n6875) );
  inv0d0 U9929 ( .I(images_bus[52]), .ZN(n6550) );
  inv0d0 U9930 ( .I(images_bus[146]), .ZN(n6778) );
  inv0d0 U9931 ( .I(images_bus[3]), .ZN(n5315) );
  inv0d0 U9932 ( .I(images_bus[392]), .ZN(n7127) );
  inv0d0 U9933 ( .I(images_bus[95]), .ZN(n6138) );
  inv0d0 U9934 ( .I(images_bus[360]), .ZN(n7133) );
  inv0d0 U9936 ( .I(images_bus[362]), .ZN(n6838) );
  inv0d0 U9937 ( .I(images_bus[124]), .ZN(n6488) );
  inv0d0 U9938 ( .I(images_bus[54]), .ZN(n6270) );
  inv0d0 U9939 ( .I(images_bus[348]), .ZN(n6445) );
  inv0d0 U9940 ( .I(images_bus[118]), .ZN(n6267) );
  inv0d0 U9941 ( .I(images_bus[426]), .ZN(n6826) );
  inv0d0 U9947 ( .I(images_bus[383]), .ZN(n6089) );
  inv0d0 U9948 ( .I(images_bus[498]), .ZN(n6723) );
  inv0d0 U9949 ( .I(images_bus[8]), .ZN(n7184) );
  inv0d0 U9950 ( .I(images_bus[246]), .ZN(n6246) );
  inv0d0 U9952 ( .I(images_bus[46]), .ZN(n6348) );
  inv0d0 U9953 ( .I(images_bus[66]), .ZN(n6953) );
  inv0d0 U9954 ( .I(images_bus[62]), .ZN(n6200) );
  inv0d0 U9955 ( .I(images_bus[318]), .ZN(n6170) );
  inv0d0 U9957 ( .I(images_bus[172]), .ZN(n6572) );
  inv0d0 U9958 ( .I(images_bus[422]), .ZN(n6360) );
  inv0d0 U9960 ( .I(images_bus[372]), .ZN(n6525) );
  inv0d0 U9961 ( .I(images_bus[100]), .ZN(n6639) );
  inv0d0 U9962 ( .I(images_bus[30]), .ZN(n6207) );
  inv0d0 U9963 ( .I(images_bus[506]), .ZN(n6654) );
  inv0d0 U9964 ( .I(images_bus[26]), .ZN(n6707) );
  inv0d0 U9965 ( .I(images_bus[23]), .ZN(n5864) );
  inv0d0 U9966 ( .I(images_bus[466]), .ZN(n6731) );
  inv0d0 U9967 ( .I(images_bus[60]), .ZN(n6502) );
  inv0d0 U9968 ( .I(images_bus[212]), .ZN(n6540) );
  inv0d0 U9969 ( .I(images_bus[273]), .ZN(n5540) );
  inv0d0 U9970 ( .I(images_bus[330]), .ZN(n6840) );
  inv0d0 U9971 ( .I(images_bus[394]), .ZN(n6837) );
  inv0d0 U9972 ( .I(images_bus[509]), .ZN(n2809) );
  inv0d0 U9973 ( .I(images_bus[238]), .ZN(n6310) );
  inv0d0 U9974 ( .I(images_bus[110]), .ZN(n6344) );
  inv0d0 U9976 ( .I(images_bus[261]), .ZN(n4689) );
  inv0d0 U9977 ( .I(images_bus[5]), .ZN(n4871) );
  inv0d0 U9978 ( .I(images_bus[186]), .ZN(n6683) );
  inv0d0 U9979 ( .I(images_bus[250]), .ZN(n6677) );
  inv0d0 U9980 ( .I(images_bus[302]), .ZN(n6303) );
  inv0d0 U9981 ( .I(images_bus[78]), .ZN(n6345) );
  inv0d0 U9982 ( .I(images_bus[33]), .ZN(n5782) );
  inv0d0 U9983 ( .I(images_bus[306]), .ZN(n6752) );
  nd03d1 U9986 ( .A1(n4309), .A2(images_bus[268]), .A3(n5413), .ZN(n7407) );
  nr02d1 U9987 ( .A1(n11124), .A2(n12125), .ZN(n11192) );
  nd03d1 U9989 ( .A1(images_bus[195]), .A2(images_bus[193]), .A3(
        images_bus[194]), .ZN(n6626) );
  inv0d0 U9992 ( .I(n9290), .ZN(n3491) );
  inv0d0 U9993 ( .I(n8272), .ZN(n4125) );
  inv0d0 U9994 ( .I(n11924), .ZN(n2880) );
  nr02d1 U9995 ( .A1(n6557), .A2(n8728), .ZN(n8727) );
  inv0d0 U9998 ( .I(n10366), .ZN(n2958) );
  nd02d1 U9999 ( .A1(n7919), .A2(n6084), .ZN(n11821) );
  inv0d0 U10000 ( .I(N13682), .ZN(n7606) );
  inv0d0 U10001 ( .I(n6609), .ZN(n3518) );
  nd03d1 U10003 ( .A1(images_bus[37]), .A2(n4286), .A3(images_bus[38]), .ZN(
        n8887) );
  nr02d1 U10004 ( .A1(n10915), .A2(n12138), .ZN(n11232) );
  nr02d1 U10005 ( .A1(n3664), .A2(n12121), .ZN(n11255) );
  nd02d1 U10006 ( .A1(n5833), .A2(images_bus[313]), .ZN(n12020) );
  nd02d1 U10007 ( .A1(n10548), .A2(n6699), .ZN(n11282) );
  nr02d1 U10008 ( .A1(n6701), .A2(n4293), .ZN(n11291) );
  nr02d1 U10010 ( .A1(n12139), .A2(n3137), .ZN(n11223) );
  nr02d1 U10011 ( .A1(n7136), .A2(n10868), .ZN(n11235) );
  nr02d1 U10012 ( .A1(n6356), .A2(n11131), .ZN(n11188) );
  nr02d1 U10013 ( .A1(n7104), .A2(n4140), .ZN(n11284) );
  nd03d1 U10014 ( .A1(n3249), .A2(n5730), .A3(n3250), .ZN(n11783) );
  nd02d1 U10015 ( .A1(n3761), .A2(n10722), .ZN(n11599) );
  nr02d1 U10017 ( .A1(n8752), .A2(n12129), .ZN(n4804) );
  nd02d1 U10018 ( .A1(n10571), .A2(n6795), .ZN(n11280) );
  nd02d1 U10019 ( .A1(n6179), .A2(n10667), .ZN(n11263) );
  nd02d1 U10020 ( .A1(n6328), .A2(n11268), .ZN(n11267) );
  aoim22d1 U10021 ( .A1(n8967), .A2(n11371), .B1(n8974), .B2(images_bus[55]), 
        .Z(n11370) );
  nr02d1 U10022 ( .A1(n10688), .A2(n12155), .ZN(n6955) );
  inv0d0 U10023 ( .I(n10292), .ZN(n2820) );
  aoim22d1 U10025 ( .A1(n10294), .A2(n2860), .B1(n10295), .B2(n10296), .Z(
        n10293) );
  nd02d1 U10026 ( .A1(n3014), .A2(n10216), .ZN(n10215) );
  nr02d1 U10027 ( .A1(n6181), .A2(n7401), .ZN(n7082) );
  inv0d0 U10029 ( .I(n8919), .ZN(n4552) );
  inv0d0 U10030 ( .I(n8921), .ZN(n4524) );
  nd02d1 U10031 ( .A1(n3168), .A2(images_bus[381]), .ZN(n6362) );
  nd02d1 U10032 ( .A1(images_bus[132]), .A2(n3988), .ZN(n11276) );
  nd02d1 U10033 ( .A1(images_bus[454]), .A2(n11083), .ZN(n11205) );
  nd02d1 U10034 ( .A1(images_bus[76]), .A2(n10530), .ZN(n11285) );
  nd02d1 U10035 ( .A1(images_bus[48]), .A2(n10498), .ZN(n11292) );
  nd02d1 U10036 ( .A1(images_bus[496]), .A2(n2815), .ZN(n11185) );
  nd02d1 U10037 ( .A1(images_bus[244]), .A2(n3660), .ZN(n11254) );
  inv0d0 U10038 ( .I(n7094), .ZN(n3455) );
  nr02d1 U10039 ( .A1(n6390), .A2(n12170), .ZN(n5765) );
  nd02d1 U10040 ( .A1(n6952), .A2(images_bus[207]), .ZN(n6949) );
  inv0d0 U10043 ( .I(n7416), .ZN(n3891) );
  inv0d0 U10044 ( .I(n4424), .ZN(n3916) );
  inv0d0 U10045 ( .I(n2258), .ZN(n2261) );
  nd02d1 U10046 ( .A1(images_bus[426]), .A2(n6460), .ZN(n7938) );
  nd02d1 U10047 ( .A1(images_bus[156]), .A2(images_bus[155]), .ZN(n5112) );
  nd02d1 U10048 ( .A1(images_bus[316]), .A2(images_bus[315]), .ZN(n4993) );
  inv0d0 U10052 ( .I(n6721), .ZN(n4252) );
  inv0d0 U10053 ( .I(n10750), .ZN(n3659) );
  nd02d1 U10054 ( .A1(n7140), .A2(n7146), .ZN(n7144) );
  inv0d0 U10055 ( .I(n7039), .ZN(n3513) );
  inv0d0 U10056 ( .I(n6980), .ZN(n3621) );
  nr02d1 U10057 ( .A1(n6634), .A2(n5989), .ZN(n6633) );
  nd03d1 U10058 ( .A1(n3963), .A2(images_bus[168]), .A3(N10266), .ZN(n5144) );
  nr02d1 U10059 ( .A1(n6367), .A2(n12124), .ZN(n4968) );
  nd02d1 U10060 ( .A1(images_bus[156]), .A2(n10619), .ZN(n11270) );
  nd02d1 U10061 ( .A1(images_bus[338]), .A2(n10879), .ZN(n11234) );
  nd03d1 U10062 ( .A1(n5344), .A2(n3097), .A3(n9487), .ZN(n9485) );
  nd02d1 U10063 ( .A1(images_bus[366]), .A2(n3269), .ZN(n11226) );
  nr02d1 U10065 ( .A1(n5523), .A2(n12132), .ZN(n4975) );
  nd02d1 U10066 ( .A1(images_bus[436]), .A2(n3020), .ZN(n11211) );
  nr13d1 U10069 ( .A1(n6831), .A2(n6832), .A3(n4133), .ZN(n6828) );
  inv0d0 U10070 ( .I(n8233), .ZN(n4217) );
  inv0d0 U10071 ( .I(n8115), .ZN(n4203) );
  inv0d0 U10073 ( .I(n10736), .ZN(n2811) );
  nd02d1 U10074 ( .A1(images_bus[44]), .A2(n4295), .ZN(n11293) );
  nd03d1 U10075 ( .A1(images_bus[344]), .A2(n3342), .A3(images_bus[345]), .ZN(
        n9364) );
  nr02d1 U10076 ( .A1(n5231), .A2(n12141), .ZN(n8045) );
  aoim22d1 U10077 ( .A1(n8361), .A2(n11535), .B1(n3926), .B2(n11536), .Z(
        n11530) );
  inv0d0 U10078 ( .I(n8358), .ZN(n3925) );
  inv0d0 U10079 ( .I(n6779), .ZN(n4132) );
  inv0d0 U10080 ( .I(n7718), .ZN(n3755) );
  nd03d1 U10081 ( .A1(n4826), .A2(n9524), .A3(n8772), .ZN(n9522) );
  nd03d1 U10083 ( .A1(images_bus[182]), .A2(n9139), .A3(images_bus[183]), .ZN(
        n11552) );
  inv0d0 U10084 ( .I(n9449), .ZN(n3032) );
  inv0d0 U10085 ( .I(n9551), .ZN(n2848) );
  inv0d0 U10086 ( .I(n4517), .ZN(n3440) );
  inv0d0 U10087 ( .I(n4906), .ZN(n2887) );
  nr13d1 U10088 ( .A1(n6143), .A2(n9259), .A3(n10786), .ZN(n10785) );
  inv0d0 U10089 ( .I(n9261), .ZN(n3544) );
  inv0d0 U10090 ( .I(n9967), .ZN(n3587) );
  nd03d1 U10091 ( .A1(n2845), .A2(n6425), .A3(n2914), .ZN(n9547) );
  inv0d0 U10092 ( .I(n10307), .ZN(n2866) );
  inv0d0 U10093 ( .I(n4391), .ZN(n4005) );
  nr02d1 U10094 ( .A1(n5669), .A2(n12128), .ZN(n8401) );
  inv0d0 U10095 ( .I(n7320), .ZN(n2928) );
  inv0d0 U10096 ( .I(n6167), .ZN(n3427) );
  nr02d1 U10097 ( .A1(n6838), .A2(n12165), .ZN(n7382) );
  inv0d0 U10098 ( .I(n10678), .ZN(n3816) );
  nr02d1 U10099 ( .A1(n6628), .A2(n12170), .ZN(n7420) );
  inv0d0 U10100 ( .I(n10608), .ZN(n3987) );
  nd02d1 U10101 ( .A1(images_bus[160]), .A2(n10624), .ZN(n11269) );
  nr02d1 U10103 ( .A1(n9968), .A2(n6174), .ZN(n10404) );
  nr02d1 U10104 ( .A1(n6747), .A2(n5825), .ZN(n7389) );
  nr02d1 U10105 ( .A1(n5418), .A2(images_bus[317]), .ZN(n7812) );
  nd02d1 U10107 ( .A1(images_bus[268]), .A2(n10774), .ZN(n11247) );
  nd02d1 U10108 ( .A1(images_bus[346]), .A2(n10898), .ZN(n11233) );
  nd02d1 U10109 ( .A1(images_bus[422]), .A2(images_bus[421]), .ZN(n4953) );
  nd02d1 U10110 ( .A1(images_bus[118]), .A2(n11279), .ZN(n11278) );
  nd02d1 U10111 ( .A1(images_bus[194]), .A2(n10671), .ZN(n11262) );
  nr02d1 U10112 ( .A1(n10240), .A2(n12156), .ZN(n8763) );
  nd02d1 U10113 ( .A1(n6737), .A2(n10936), .ZN(n11224) );
  nd03d1 U10114 ( .A1(N14386), .A2(n11833), .A3(images_bus[431]), .ZN(n5600)
         );
  nd02d1 U10115 ( .A1(images_bus[122]), .A2(images_bus[121]), .ZN(n6825) );
  inv0d0 U10116 ( .I(n10167), .ZN(n3133) );
  inv0d0 U10117 ( .I(n5821), .ZN(n4147) );
  nr02d1 U10118 ( .A1(n5398), .A2(n5636), .ZN(n6607) );
  nr02d1 U10120 ( .A1(n5831), .A2(images_bus[77]), .ZN(n8251) );
  nd02d1 U10121 ( .A1(images_bus[124]), .A2(images_bus[123]), .ZN(n6650) );
  nd02d1 U10122 ( .A1(images_bus[250]), .A2(images_bus[249]), .ZN(n7411) );
  nd03d1 U10125 ( .A1(N14034), .A2(n3224), .A3(images_bus[409]), .ZN(n8658) );
  nd02d1 U10126 ( .A1(images_bus[89]), .A2(n6699), .ZN(n7447) );
  nd02d1 U10127 ( .A1(images_bus[178]), .A2(n11266), .ZN(n11265) );
  nd03d1 U10128 ( .A1(images_bus[182]), .A2(n9139), .A3(N10476), .ZN(n6917) );
  nd03d1 U10129 ( .A1(n11857), .A2(n4635), .A3(n8041), .ZN(n11856) );
  inv0d0 U10130 ( .I(n6026), .ZN(n3898) );
  nd03d1 U10131 ( .A1(n11681), .A2(images_bus[307]), .A3(N12402), .ZN(n7090)
         );
  inv0d0 U10132 ( .I(n8832), .ZN(n2846) );
  inv0d0 U10133 ( .I(n2244), .ZN(n2247) );
  nd03d1 U10134 ( .A1(n4171), .A2(n4163), .A3(n4166), .ZN(n6767) );
  nd02d1 U10135 ( .A1(images_bus[248]), .A2(images_bus[247]), .ZN(n5330) );
  inv0d0 U10136 ( .I(n6444), .ZN(n3130) );
  inv0d0 U10137 ( .I(n5103), .ZN(n4041) );
  nd03d1 U10138 ( .A1(n9346), .A2(n10884), .A3(n3404), .ZN(n10876) );
  nd03d1 U10139 ( .A1(images_bus[204]), .A2(n9167), .A3(N10806), .ZN(n11259)
         );
  nd02d1 U10140 ( .A1(images_bus[409]), .A2(n6659), .ZN(n5709) );
  nd02d1 U10141 ( .A1(images_bus[205]), .A2(n6324), .ZN(n5218) );
  nd03d1 U10142 ( .A1(n9076), .A2(images_bus[119]), .A3(N9540), .ZN(n5030) );
  nd02d1 U10143 ( .A1(images_bus[418]), .A2(images_bus[417]), .ZN(n4955) );
  inv0d0 U10144 ( .I(n6797), .ZN(n4109) );
  inv0d0 U10145 ( .I(n6454), .ZN(n3124) );
  inv0d0 U10148 ( .I(n10346), .ZN(n2901) );
  nd02d1 U10149 ( .A1(images_bus[498]), .A2(images_bus[497]), .ZN(n4919) );
  inv0d0 U10150 ( .I(n5030), .ZN(n4088) );
  nd03d1 U10151 ( .A1(n6561), .A2(images_bus[438]), .A3(n6477), .ZN(n6483) );
  nd02d1 U10152 ( .A1(images_bus[167]), .A2(images_bus[168]), .ZN(n5139) );
  nd03d1 U10153 ( .A1(N14706), .A2(n3008), .A3(images_bus[451]), .ZN(n4791) );
  inv0d0 U10154 ( .I(n8984), .ZN(n4282) );
  nd02d1 U10155 ( .A1(images_bus[380]), .A2(images_bus[379]), .ZN(n4969) );
  nr02d1 U10156 ( .A1(n6685), .A2(n12120), .ZN(n6688) );
  nr02d1 U10157 ( .A1(n8112), .A2(n8111), .ZN(n7535) );
  nd02d1 U10158 ( .A1(images_bus[231]), .A2(n7153), .ZN(n5296) );
  aoim22d1 U10159 ( .A1(n4442), .A2(n9238), .B1(n9242), .B2(n9243), .Z(n9241)
         );
  nd02d1 U10160 ( .A1(images_bus[366]), .A2(images_bus[365]), .ZN(n6318) );
  nr02d1 U10161 ( .A1(n6992), .A2(n8437), .ZN(n8444) );
  nd02d1 U10162 ( .A1(n3161), .A2(images_bus[383]), .ZN(n4970) );
  inv0d0 U10163 ( .I(n5236), .ZN(n3852) );
  nd02d1 U10164 ( .A1(images_bus[348]), .A2(images_bus[347]), .ZN(n4982) );
  nd02d1 U10165 ( .A1(images_bus[217]), .A2(n6682), .ZN(n5757) );
  nd03d1 U10166 ( .A1(n8197), .A2(images_bus[45]), .A3(N8523), .ZN(n6713) );
  nd03d1 U10167 ( .A1(images_bus[494]), .A2(n2882), .A3(N15394), .ZN(n8810) );
  nd02d1 U10168 ( .A1(images_bus[188]), .A2(n4958), .ZN(n5769) );
  nd02d1 U10169 ( .A1(images_bus[126]), .A2(images_bus[125]), .ZN(n6649) );
  nr02d1 U10170 ( .A1(n5607), .A2(n12129), .ZN(n7317) );
  nd03d1 U10171 ( .A1(N14114), .A2(n6430), .A3(images_bus[414]), .ZN(n8679) );
  nd02d1 U10172 ( .A1(images_bus[310]), .A2(images_bus[309]), .ZN(n7396) );
  nd02d1 U10173 ( .A1(images_bus[110]), .A2(images_bus[109]), .ZN(n7442) );
  inv0d0 U10174 ( .I(n8206), .ZN(n2793) );
  nd02d1 U10175 ( .A1(images_bus[182]), .A2(images_bus[181]), .ZN(n5774) );
  nd03d1 U10176 ( .A1(images_bus[204]), .A2(n9167), .A3(images_bus[205]), .ZN(
        n10688) );
  nd02d1 U10177 ( .A1(images_bus[400]), .A2(images_bus[399]), .ZN(n4963) );
  nd03d1 U10178 ( .A1(n9104), .A2(images_bus[141]), .A3(N9861), .ZN(n5967) );
  aoim22d1 U10179 ( .A1(n7058), .A2(n3471), .B1(n5388), .B2(images_bus[293]), 
        .Z(n7054) );
  aoim22d1 U10180 ( .A1(n5789), .A2(n6712), .B1(n6713), .B2(n6714), .Z(n6708)
         );
  nd02d1 U10182 ( .A1(images_bus[419]), .A2(n6599), .ZN(n7366) );
  nr02d1 U10183 ( .A1(n9836), .A2(images_bus[147]), .ZN(n5090) );
  nd02d1 U10184 ( .A1(images_bus[373]), .A2(n8601), .ZN(n5504) );
  nd03d1 U10186 ( .A1(images_bus[311]), .A2(n10837), .A3(N12466), .ZN(n9312)
         );
  nd03d1 U10187 ( .A1(N15122), .A2(n11898), .A3(images_bus[477]), .ZN(n9542)
         );
  nd03d1 U10188 ( .A1(n10402), .A2(images_bus[259]), .A3(N11634), .ZN(n10762)
         );
  nd03d1 U10189 ( .A1(n12059), .A2(images_bus[189]), .A3(N10581), .ZN(n5193)
         );
  nd02d1 U10190 ( .A1(images_bus[289]), .A2(n6922), .ZN(n4483) );
  nd02d1 U10191 ( .A1(images_bus[404]), .A2(images_bus[403]), .ZN(n7375) );
  inv0d0 U10192 ( .I(n9214), .ZN(n3717) );
  inv0d0 U10193 ( .I(n5064), .ZN(n2806) );
  nd03d1 U10194 ( .A1(N14834), .A2(n4804), .A3(images_bus[459]), .ZN(n7319) );
  nr02d1 U10195 ( .A1(n5334), .A2(images_bus[249]), .ZN(n7740) );
  nd03d1 U10196 ( .A1(n4305), .A2(images_bus[375]), .A3(n8604), .ZN(n8608) );
  nd02d1 U10198 ( .A1(images_bus[384]), .A2(n11779), .ZN(n7215) );
  nd02d1 U10199 ( .A1(images_bus[172]), .A2(images_bus[171]), .ZN(n7430) );
  nd02d1 U10200 ( .A1(images_bus[238]), .A2(images_bus[237]), .ZN(n5308) );
  nd03d1 U10201 ( .A1(images_bus[346]), .A2(n12004), .A3(N13026), .ZN(n8570)
         );
  nd03d1 U10203 ( .A1(n3879), .A2(n7685), .A3(images_bus[201]), .ZN(n5209) );
  nd02d1 U10205 ( .A1(images_bus[186]), .A2(images_bus[185]), .ZN(n6631) );
  nd02d1 U10206 ( .A1(images_bus[457]), .A2(n7311), .ZN(n8752) );
  nd02d1 U10207 ( .A1(images_bus[210]), .A2(images_bus[209]), .ZN(n5234) );
  nr02d1 U10209 ( .A1(n5242), .A2(n12139), .ZN(n4645) );
  an03d1 U10210 ( .A1(n1344), .A2(n11622), .A3(images_bus[254]), .Z(n5348) );
  nd02d1 U10211 ( .A1(images_bus[108]), .A2(n5911), .ZN(n8290) );
  nd02d1 U10212 ( .A1(images_bus[326]), .A2(images_bus[325]), .ZN(n4990) );
  nd03d1 U10213 ( .A1(images_bus[86]), .A2(n11286), .A3(N9078), .ZN(n5859) );
  nd02d1 U10214 ( .A1(images_bus[368]), .A2(images_bus[367]), .ZN(n6597) );
  nd03d1 U10215 ( .A1(n2886), .A2(images_bus[497]), .A3(N15442), .ZN(n11156)
         );
  nd02d1 U10216 ( .A1(images_bus[60]), .A2(images_bus[59]), .ZN(n8222) );
  nr02d1 U10217 ( .A1(n8081), .A2(n7714), .ZN(n8080) );
  nd03d1 U10218 ( .A1(n4079), .A2(images_bus[109]), .A3(N9400), .ZN(n5917) );
  nd03d1 U10219 ( .A1(images_bus[484]), .A2(n10288), .A3(images_bus[485]), 
        .ZN(n11130) );
  nd02d1 U10221 ( .A1(images_bus[334]), .A2(n12012), .ZN(n8563) );
  nd03d1 U10222 ( .A1(n4055), .A2(images_bus[132]), .A3(N9726), .ZN(n9638) );
  nd03d1 U10223 ( .A1(images_bus[15]), .A2(n8147), .A3(images_bus[16]), .ZN(
        n10452) );
  nd02d1 U10224 ( .A1(images_bus[158]), .A2(images_bus[157]), .ZN(n7645) );
  nd03d1 U10226 ( .A1(n4113), .A2(images_bus[101]), .A3(N9288), .ZN(n9050) );
  inv0d0 U10229 ( .I(n6876), .ZN(n3900) );
  nd02d1 U10230 ( .A1(n5771), .A2(images_bus[130]), .ZN(n5053) );
  nd02d1 U10231 ( .A1(n2934), .A2(images_bus[448]), .ZN(n4942) );
  nd03d1 U10232 ( .A1(images_bus[474]), .A2(n2980), .A3(N15074), .ZN(n8781) );
  nd02d1 U10233 ( .A1(images_bus[328]), .A2(images_bus[327]), .ZN(n4989) );
  nd02d1 U10234 ( .A1(finish_flag), .A2(N8001), .ZN(n5008) );
  inv0d0 U10235 ( .I(n6620), .ZN(n3576) );
  nd02d1 U10236 ( .A1(images_bus[189]), .A2(n6179), .ZN(n6935) );
  nd02d1 U10237 ( .A1(images_bus[463]), .A2(n8763), .ZN(n9525) );
  inv0d0 U10240 ( .I(n9720), .ZN(n4225) );
  nd02d1 U10243 ( .A1(images_bus[464]), .A2(n2993), .ZN(n10368) );
  nd02d1 U10244 ( .A1(images_bus[296]), .A2(images_bus[295]), .ZN(n5398) );
  nd02d1 U10247 ( .A1(images_bus[496]), .A2(n11931), .ZN(n8813) );
  nr02d1 U10248 ( .A1(n7583), .A2(n12131), .ZN(n10568) );
  nd03d1 U10249 ( .A1(images_bus[84]), .A2(n11416), .A3(N9050), .ZN(n6768) );
  nd03d1 U10255 ( .A1(n5904), .A2(n11833), .A3(images_bus[433]), .ZN(n7955) );
  nd03d1 U10256 ( .A1(images_bus[293]), .A2(n5384), .A3(N12178), .ZN(n5392) );
  nd03d1 U10257 ( .A1(n4439), .A2(n3461), .A3(images_bus[303]), .ZN(n6183) );
  inv0d0 U10258 ( .I(n6326), .ZN(n3311) );
  aoim22d1 U10259 ( .A1(n6331), .A2(n7196), .B1(n5500), .B2(images_bus[375]), 
        .Z(n7195) );
  nd03d1 U10260 ( .A1(images_bus[404]), .A2(n11220), .A3(N13954), .ZN(n6409)
         );
  nd03d1 U10261 ( .A1(images_bus[104]), .A2(n8282), .A3(N9330), .ZN(n5905) );
  nd02d1 U10262 ( .A1(images_bus[225]), .A2(n6931), .ZN(n5755) );
  nd03d1 U10263 ( .A1(N14290), .A2(n8691), .A3(images_bus[425]), .ZN(n9471) );
  inv0d0 U10264 ( .I(n1623), .ZN(n1626) );
  inv0d0 U10265 ( .I(n9964), .ZN(n3586) );
  nd03d1 U10266 ( .A1(N14002), .A2(n3234), .A3(images_bus[407]), .ZN(n6421) );
  nd02d1 U10267 ( .A1(images_bus[113]), .A2(n6795), .ZN(n5926) );
  inv0d0 U10269 ( .I(n7570), .ZN(n4130) );
  nd02d1 U10270 ( .A1(images_bus[82]), .A2(images_bus[81]), .ZN(n6662) );
  nd02d1 U10271 ( .A1(images_bus[222]), .A2(images_bus[221]), .ZN(n7711) );
  nd02d1 U10272 ( .A1(images_bus[234]), .A2(images_bus[233]), .ZN(n7413) );
  nr02d1 U10273 ( .A1(n5388), .A2(images_bus[293]), .ZN(n4997) );
  nd03d1 U10274 ( .A1(images_bus[274]), .A2(n5362), .A3(N11874), .ZN(n5358) );
  inv0d0 U10275 ( .I(n1998), .ZN(n1999) );
  nd02d1 U10277 ( .A1(images_bus[214]), .A2(images_bus[213]), .ZN(n7704) );
  nd03d1 U10278 ( .A1(n2902), .A2(images_bus[507]), .A3(N15602), .ZN(n11182)
         );
  nd02d1 U10279 ( .A1(images_bus[242]), .A2(images_bus[241]), .ZN(n6106) );
  nd03d1 U10280 ( .A1(n4308), .A2(images_bus[311]), .A3(n9302), .ZN(n9311) );
  nr02d1 U10281 ( .A1(n9227), .A2(images_bus[247]), .ZN(n5332) );
  inv0d0 U10282 ( .I(n8837), .ZN(n3237) );
  nd03d1 U10284 ( .A1(images_bus[491]), .A2(n11932), .A3(N15346), .ZN(n8828)
         );
  inv0d0 U10288 ( .I(n8144), .ZN(n4776) );
  nr02d1 U10289 ( .A1(n5585), .A2(n12130), .ZN(n8118) );
  nr02d1 U10290 ( .A1(n4321), .A2(n12143), .ZN(n9072) );
  nr02d1 U10291 ( .A1(n6641), .A2(n11384), .ZN(n12069) );
  nd02d1 U10292 ( .A1(images_bus[113]), .A2(n12065), .ZN(n7583) );
  nd02d1 U10293 ( .A1(images_bus[240]), .A2(images_bus[239]), .ZN(n6619) );
  nr02d1 U10294 ( .A1(images_bus[423]), .A2(n9469), .ZN(n9467) );
  nd02d1 U10295 ( .A1(images_bus[33]), .A2(images_bus[32]), .ZN(n6685) );
  inv0d0 U10296 ( .I(N8044), .ZN(n7586) );
  inv0d0 U10297 ( .I(n9604), .ZN(n3217) );
  nd03d1 U10298 ( .A1(images_bus[207]), .A2(n6955), .A3(N10851), .ZN(n5225) );
  nd02d1 U10299 ( .A1(images_bus[63]), .A2(n8884), .ZN(n7452) );
  nd03d1 U10300 ( .A1(n8988), .A2(images_bus[61]), .A3(N8731), .ZN(n8992) );
  nd02d1 U10301 ( .A1(images_bus[156]), .A2(n4045), .ZN(n5109) );
  nd03d1 U10302 ( .A1(n5870), .A2(images_bus[21]), .A3(n8921), .ZN(n8926) );
  nd03d1 U10303 ( .A1(images_bus[166]), .A2(n3964), .A3(images_bus[167]), .ZN(
        n5994) );
  inv0d0 U10304 ( .I(n11411), .ZN(n4143) );
  nd02d1 U10306 ( .A1(images_bus[423]), .A2(n3126), .ZN(n11828) );
  nd03d1 U10308 ( .A1(images_bus[276]), .A2(n3559), .A3(N11906), .ZN(n9259) );
  nd03d1 U10309 ( .A1(images_bus[502]), .A2(n2892), .A3(N15522), .ZN(n9578) );
  nd02d1 U10310 ( .A1(images_bus[318]), .A2(images_bus[317]), .ZN(n4526) );
  inv0d0 U10311 ( .I(n9563), .ZN(n2881) );
  nd03d1 U10312 ( .A1(n3467), .A2(images_bus[297]), .A3(N12242), .ZN(n10823)
         );
  inv0d0 U10313 ( .I(n9394), .ZN(n3287) );
  inv0d0 U10314 ( .I(n5739), .ZN(n3511) );
  inv0d0 U10315 ( .I(n5429), .ZN(n3363) );
  nd02d1 U10316 ( .A1(images_bus[46]), .A2(images_bus[45]), .ZN(n8204) );
  nd02d1 U10317 ( .A1(images_bus[71]), .A2(images_bus[70]), .ZN(n6748) );
  inv0d0 U10318 ( .I(n5132), .ZN(n3919) );
  nd02d1 U10320 ( .A1(images_bus[108]), .A2(images_bus[107]), .ZN(n5918) );
  inv0d0 U10321 ( .I(n4539), .ZN(n3417) );
  nd02d1 U10322 ( .A1(images_bus[431]), .A2(n7062), .ZN(n5702) );
  nd02d1 U10323 ( .A1(images_bus[507]), .A2(n6423), .ZN(n8020) );
  nd03d1 U10324 ( .A1(n6271), .A2(images_bus[350]), .A3(N13090), .ZN(n10086)
         );
  nd03d1 U10325 ( .A1(n10657), .A2(images_bus[185]), .A3(N10521), .ZN(n6927)
         );
  nd02d1 U10326 ( .A1(images_bus[170]), .A2(images_bus[169]), .ZN(n7433) );
  nd03d1 U10327 ( .A1(n8774), .A2(n5798), .A3(n9539), .ZN(n9537) );
  nd02d1 U10328 ( .A1(images_bus[493]), .A2(n2910), .ZN(n11187) );
  nd02d1 U10329 ( .A1(images_bus[118]), .A2(images_bus[117]), .ZN(n5936) );
  inv0d0 U10331 ( .I(n10146), .ZN(n3139) );
  nd02d1 U10332 ( .A1(images_bus[154]), .A2(images_bus[153]), .ZN(n7640) );
  nd02d1 U10334 ( .A1(images_bus[307]), .A2(n6531), .ZN(n7400) );
  nd03d1 U10335 ( .A1(n4269), .A2(images_bus[51]), .A3(N8601), .ZN(n8214) );
  nd03d1 U10336 ( .A1(N15154), .A2(n2849), .A3(images_bus[479]), .ZN(n8796) );
  nr02d1 U10337 ( .A1(n6363), .A2(n12124), .ZN(n11997) );
  nd02d1 U10338 ( .A1(images_bus[43]), .A2(images_bus[42]), .ZN(n7457) );
  nd02d1 U10339 ( .A1(images_bus[492]), .A2(images_bus[491]), .ZN(n4924) );
  nd03d1 U10342 ( .A1(images_bus[166]), .A2(n3964), .A3(N10236), .ZN(n5135) );
  nd03d1 U10343 ( .A1(n2908), .A2(n4297), .A3(images_bus[500]), .ZN(n9574) );
  nd03d1 U10344 ( .A1(n3804), .A2(images_bus[237]), .A3(N11301), .ZN(n8445) );
  nr02d1 U10345 ( .A1(n4306), .A2(n12157), .ZN(n5723) );
  nd02d1 U10346 ( .A1(images_bus[194]), .A2(n5756), .ZN(n5766) );
  nd02d1 U10347 ( .A1(images_bus[309]), .A2(n11679), .ZN(n9304) );
  nd03d1 U10348 ( .A1(n4169), .A2(images_bus[89]), .A3(N9120), .ZN(n5866) );
  nd03d1 U10349 ( .A1(n5783), .A2(images_bus[152]), .A3(n3993), .ZN(n11508) );
  nd03d1 U10350 ( .A1(images_bus[129]), .A2(n11473), .A3(N9681), .ZN(n5948) );
  inv0d0 U10351 ( .I(n8157), .ZN(n4338) );
  nd02d1 U10352 ( .A1(images_bus[220]), .A2(images_bus[219]), .ZN(n8082) );
  nd03d1 U10353 ( .A1(images_bus[317]), .A2(n9319), .A3(N12562), .ZN(n10850)
         );
  nr02d1 U10354 ( .A1(n7115), .A2(n12166), .ZN(n9586) );
  nd02d1 U10355 ( .A1(images_bus[184]), .A2(images_bus[183]), .ZN(n6921) );
  nd03d1 U10356 ( .A1(images_bus[496]), .A2(n5124), .A3(images_bus[495]), .ZN(
        n11959) );
  nr02d1 U10357 ( .A1(n7381), .A2(images_bus[363]), .ZN(n6306) );
  nd03d1 U10358 ( .A1(n3013), .A2(images_bus[444]), .A3(n6494), .ZN(n6509) );
  nd03d1 U10359 ( .A1(n5770), .A2(images_bus[192]), .A3(N10626), .ZN(n6014) );
  nd02d1 U10360 ( .A1(n8174), .A2(images_bus[29]), .ZN(n9691) );
  nr02d1 U10361 ( .A1(n10555), .A2(images_bus[99]), .ZN(n6783) );
  nd02d1 U10362 ( .A1(images_bus[91]), .A2(n6496), .ZN(n8107) );
  nd02d1 U10363 ( .A1(images_bus[66]), .A2(n5779), .ZN(n5807) );
  nd02d1 U10364 ( .A1(images_bus[289]), .A2(n4484), .ZN(n8510) );
  nd02d1 U10365 ( .A1(images_bus[442]), .A2(n5354), .ZN(n6554) );
  nd03d1 U10366 ( .A1(n4964), .A2(images_bus[396]), .A3(n7886), .ZN(n7894) );
  nr02d1 U10367 ( .A1(n12167), .A2(n3097), .ZN(n6559) );
  nr02d1 U10369 ( .A1(n9687), .A2(images_bus[27]), .ZN(n8168) );
  nd03d1 U10370 ( .A1(n4365), .A2(images_bus[22]), .A3(N8234), .ZN(n9679) );
  nd03d1 U10372 ( .A1(n4330), .A2(images_bus[55]), .A3(n5465), .ZN(n6740) );
  nd03d1 U10373 ( .A1(N14994), .A2(n10257), .A3(images_bus[469]), .ZN(n10361)
         );
  nd02d1 U10374 ( .A1(images_bus[212]), .A2(images_bus[211]), .ZN(n8863) );
  nd02d1 U10375 ( .A1(n2935), .A2(images_bus[447]), .ZN(n8033) );
  nd02d1 U10376 ( .A1(images_bus[115]), .A2(n10568), .ZN(n6812) );
  nd03d1 U10378 ( .A1(n11968), .A2(images_bus[472]), .A3(N15042), .ZN(n11196)
         );
  nd02d1 U10379 ( .A1(images_bus[372]), .A2(images_bus[371]), .ZN(n5716) );
  nd03d1 U10380 ( .A1(n4964), .A2(images_bus[396]), .A3(n6384), .ZN(n6399) );
  nd02d1 U10381 ( .A1(images_bus[394]), .A2(images_bus[393]), .ZN(n6591) );
  nd02d1 U10382 ( .A1(images_bus[377]), .A2(n6664), .ZN(n6595) );
  nd02d1 U10383 ( .A1(images_bus[106]), .A2(images_bus[105]), .ZN(n7443) );
  nd02d1 U10384 ( .A1(images_bus[314]), .A2(images_bus[313]), .ZN(n6604) );
  nd03d1 U10385 ( .A1(images_bus[119]), .A2(n4322), .A3(n8300), .ZN(n8302) );
  nd02d1 U10386 ( .A1(images_bus[298]), .A2(images_bus[297]), .ZN(n8518) );
  nd03d1 U10387 ( .A1(n6247), .A2(images_bus[340]), .A3(images_bus[341]), .ZN(
        n5455) );
  nd03d1 U10388 ( .A1(images_bus[159]), .A2(images_bus[158]), .A3(n6865), .ZN(
        n6870) );
  nd03d1 U10389 ( .A1(images_bus[486]), .A2(n2864), .A3(N15266), .ZN(n10296)
         );
  nd02d1 U10390 ( .A1(images_bus[178]), .A2(n6910), .ZN(n8373) );
  nd03d1 U10391 ( .A1(images_bus[317]), .A2(n9319), .A3(images_bus[318]), .ZN(
        n11689) );
  nd03d1 U10392 ( .A1(N14930), .A2(n2967), .A3(images_bus[465]), .ZN(n9597) );
  nd02d1 U10393 ( .A1(images_bus[137]), .A2(n6871), .ZN(n7436) );
  nd02d1 U10394 ( .A1(images_bus[494]), .A2(images_bus[493]), .ZN(n8815) );
  nd02d1 U10396 ( .A1(images_bus[12]), .A2(n4827), .ZN(n10445) );
  nd03d1 U10397 ( .A1(images_bus[176]), .A2(images_bus[175]), .A3(n6905), .ZN(
        n6907) );
  nd02d1 U10400 ( .A1(images_bus[293]), .A2(n6383), .ZN(n6608) );
  nd02d1 U10401 ( .A1(images_bus[376]), .A2(images_bus[375]), .ZN(n6346) );
  nd02d1 U10402 ( .A1(images_bus[364]), .A2(images_bus[363]), .ZN(n4611) );
  nd02d1 U10403 ( .A1(images_bus[173]), .A2(n6328), .ZN(n7429) );
  aoim22d1 U10405 ( .A1(n8306), .A2(n8307), .B1(n5951), .B2(n8308), .Z(n8305)
         );
  nr02d1 U10406 ( .A1(n3017), .A2(images_bus[445]), .ZN(n8736) );
  nd03d1 U10407 ( .A1(images_bus[136]), .A2(images_bus[135]), .A3(n5058), .ZN(
        n5062) );
  nd02d1 U10408 ( .A1(images_bus[23]), .A2(images_bus[22]), .ZN(n7481) );
  nd03d1 U10409 ( .A1(n8045), .A2(n3008), .A3(images_bus[453]), .ZN(n11857) );
  nd03d1 U10410 ( .A1(images_bus[139]), .A2(n4024), .A3(N9831), .ZN(n8323) );
  nd03d1 U10411 ( .A1(images_bus[404]), .A2(n11220), .A3(images_bus[405]), 
        .ZN(n8644) );
  nr02d1 U10412 ( .A1(n9889), .A2(n12168), .ZN(n9887) );
  nd02d1 U10414 ( .A1(images_bus[338]), .A2(n12007), .ZN(n11716) );
  nd03d1 U10415 ( .A1(images_bus[484]), .A2(n10288), .A3(N15234), .ZN(n11194)
         );
  nd02d1 U10416 ( .A1(images_bus[67]), .A2(n4190), .ZN(n5809) );
  nr02d1 U10418 ( .A1(n8570), .A2(images_bus[347]), .ZN(n8575) );
  nd03d1 U10419 ( .A1(images_bus[222]), .A2(n3810), .A3(N11076), .ZN(n5270) );
  nd03d1 U10420 ( .A1(N13490), .A2(n6333), .A3(images_bus[375]), .ZN(n10952)
         );
  nr02d1 U10421 ( .A1(n2998), .A2(images_bus[461]), .ZN(n8760) );
  nd03d1 U10423 ( .A1(n3266), .A2(images_bus[352]), .A3(n11731), .ZN(n11733)
         );
  nd03d1 U10424 ( .A1(images_bus[96]), .A2(n8272), .A3(n5890), .ZN(n8275) );
  nd03d1 U10425 ( .A1(images_bus[96]), .A2(n8103), .A3(n5890), .ZN(n7570) );
  nd03d1 U10426 ( .A1(n7420), .A2(images_bus[195]), .A3(n8389), .ZN(n8393) );
  nd03d1 U10427 ( .A1(n5970), .A2(images_bus[143]), .A3(n8324), .ZN(n8328) );
  nd02d1 U10428 ( .A1(images_bus[357]), .A2(n7160), .ZN(n9379) );
  nd02d1 U10429 ( .A1(images_bus[464]), .A2(images_bus[463]), .ZN(n4820) );
  nd03d1 U10430 ( .A1(n3266), .A2(images_bus[352]), .A3(n4573), .ZN(n4581) );
  nd02d1 U10431 ( .A1(images_bus[488]), .A2(images_bus[487]), .ZN(n11960) );
  nd02d1 U10432 ( .A1(n3009), .A2(images_bus[450]), .ZN(n9501) );
  nr02d1 U10433 ( .A1(n10259), .A2(n12147), .ZN(n10363) );
  nr02d1 U10434 ( .A1(n4890), .A2(n12151), .ZN(n7999) );
  nd03d1 U10435 ( .A1(N11970), .A2(n12032), .A3(images_bus[280]), .ZN(n11244)
         );
  nr02d1 U10436 ( .A1(n10883), .A2(images_bus[337]), .ZN(n6241) );
  nd03d1 U10437 ( .A1(images_bus[199]), .A2(n5765), .A3(n9154), .ZN(n9628) );
  nd03d1 U10438 ( .A1(images_bus[266]), .A2(n9977), .A3(N11746), .ZN(n7028) );
  inv0d0 U10439 ( .I(reset), .ZN(n7567) );
  nd03d1 U10440 ( .A1(images_bus[207]), .A2(n6955), .A3(images_bus[208]), .ZN(
        n9911) );
  inv0d0 U10441 ( .I(n5599), .ZN(n3085) );
  nd02d1 U10442 ( .A1(images_bus[467]), .A2(n6512), .ZN(n7985) );
  nr02d1 U10443 ( .A1(n5995), .A2(images_bus[175]), .ZN(n9875) );
  aoim22d1 U10446 ( .A1(n3947), .A2(n5176), .B1(n5177), .B2(n5178), .Z(n5175)
         );
  inv0d0 U10447 ( .I(n8477), .ZN(n3565) );
  nr02d1 U10448 ( .A1(n10090), .A2(images_bus[355]), .ZN(n7149) );
  nr02d1 U10449 ( .A1(n5976), .A2(images_bus[157]), .ZN(n9122) );
  nd03d1 U10450 ( .A1(n10257), .A2(n6212), .A3(images_bus[469]), .ZN(n7332) );
  nr02d1 U10451 ( .A1(n11362), .A2(images_bus[49]), .ZN(n6724) );
  nr02d1 U10452 ( .A1(n10828), .A2(images_bus[301]), .ZN(n8523) );
  nd03d1 U10455 ( .A1(N14610), .A2(n11854), .A3(images_bus[445]), .ZN(n8737)
         );
  nd02d1 U10456 ( .A1(images_bus[94]), .A2(images_bus[93]), .ZN(n5879) );
  inv0d0 U10457 ( .I(n8954), .ZN(n4249) );
  nd03d1 U10458 ( .A1(images_bus[175]), .A2(n9876), .A3(images_bus[176]), .ZN(
        n5167) );
  nr02d1 U10459 ( .A1(n9989), .A2(images_bus[269]), .ZN(n8484) );
  nd03d1 U10461 ( .A1(n8862), .A2(n3870), .A3(images_bus[216]), .ZN(n5256) );
  nd02d1 U10462 ( .A1(images_bus[434]), .A2(images_bus[433]), .ZN(n4947) );
  inv0d0 U10463 ( .I(N14530), .ZN(n7611) );
  inv0d0 U10464 ( .I(n5908), .ZN(n4122) );
  nd03d1 U10465 ( .A1(N14514), .A2(n3112), .A3(images_bus[439]), .ZN(n6486) );
  nd02d1 U10466 ( .A1(images_bus[353]), .A2(n6908), .ZN(n4979) );
  nd03d1 U10467 ( .A1(n4093), .A2(images_bus[121]), .A3(N9568), .ZN(n7599) );
  nd02d1 U10469 ( .A1(images_bus[150]), .A2(images_bus[149]), .ZN(n8096) );
  inv0d0 U10470 ( .I(n8244), .ZN(n4148) );
  nd03d1 U10473 ( .A1(n5725), .A2(images_bus[333]), .A3(n5448), .ZN(n5446) );
  nd03d1 U10475 ( .A1(N12530), .A2(n3445), .A3(images_bus[315]), .ZN(n5420) );
  inv0d0 U10476 ( .I(n5216), .ZN(n5665) );
  nd03d1 U10477 ( .A1(n3942), .A2(images_bus[179]), .A3(N10431), .ZN(n4394) );
  nd03d1 U10478 ( .A1(n3873), .A2(images_bus[211]), .A3(N10911), .ZN(n5246) );
  nd02d1 U10479 ( .A1(images_bus[288]), .A2(n7404), .ZN(n7051) );
  nd03d1 U10480 ( .A1(n3240), .A2(n9440), .A3(n3238), .ZN(n9435) );
  nd03d1 U10481 ( .A1(n4184), .A2(images_bus[70]), .A3(N8854), .ZN(n5816) );
  nr02d1 U10482 ( .A1(n6595), .A2(n7201), .ZN(n7203) );
  nd02d1 U10483 ( .A1(images_bus[461]), .A2(n3001), .ZN(n10240) );
  nd03d1 U10484 ( .A1(n6247), .A2(images_bus[340]), .A3(N12930), .ZN(n6253) );
  nd03d1 U10485 ( .A1(images_bus[309]), .A2(n5052), .A3(n5408), .ZN(n5411) );
  nd03d1 U10486 ( .A1(images_bus[175]), .A2(n4470), .A3(n9129), .ZN(n9136) );
  nd02d1 U10487 ( .A1(n4438), .A2(images_bus[303]), .ZN(n5733) );
  nd02d1 U10488 ( .A1(n5075), .A2(images_bus[140]), .ZN(n5072) );
  inv0d0 U10489 ( .I(n4502), .ZN(n3430) );
  nd02d1 U10490 ( .A1(images_bus[399]), .A2(n7227), .ZN(n6394) );
  nr02d1 U10491 ( .A1(n6252), .A2(images_bus[339]), .ZN(n6249) );
  nd02d1 U10492 ( .A1(images_bus[136]), .A2(n6851), .ZN(n7619) );
  nd02d1 U10493 ( .A1(images_bus[314]), .A2(n11680), .ZN(n10045) );
  nd02d1 U10494 ( .A1(n9963), .A2(images_bus[247]), .ZN(n9964) );
  nd03d1 U10495 ( .A1(N12210), .A2(n7064), .A3(images_bus[295]), .ZN(n10020)
         );
  inv0d0 U10496 ( .I(n1947), .ZN(n1950) );
  nd02d1 U10497 ( .A1(images_bus[433]), .A2(n7062), .ZN(n8720) );
  nd03d1 U10498 ( .A1(images_bus[57]), .A2(n12071), .A3(images_bus[58]), .ZN(
        n11378) );
  nd02d1 U10499 ( .A1(images_bus[416]), .A2(n11981), .ZN(n7918) );
  nd03d1 U10500 ( .A1(images_bus[324]), .A2(n4537), .A3(n3348), .ZN(n11705) );
  nd03d1 U10501 ( .A1(images_bus[17]), .A2(n4590), .A3(images_bus[18]), .ZN(
        n11325) );
  nd03d1 U10502 ( .A1(images_bus[103]), .A2(n6657), .A3(n9042), .ZN(n9048) );
  nd03d1 U10503 ( .A1(images_bus[106]), .A2(n6790), .A3(N9358), .ZN(n7578) );
  nd02d1 U10504 ( .A1(images_bus[406]), .A2(images_bus[405]), .ZN(n6415) );
  nd03d1 U10505 ( .A1(images_bus[126]), .A2(n4057), .A3(images_bus[127]), .ZN(
        n8311) );
  nd02d1 U10506 ( .A1(images_bus[392]), .A2(images_bus[391]), .ZN(n5713) );
  nd02d1 U10507 ( .A1(images_bus[411]), .A2(n6437), .ZN(n5708) );
  nd02d1 U10508 ( .A1(images_bus[360]), .A2(images_bus[359]), .ZN(n6296) );
  nd02d1 U10509 ( .A1(images_bus[236]), .A2(images_bus[235]), .ZN(n8858) );
  nd03d1 U10510 ( .A1(N15490), .A2(n2908), .A3(images_bus[500]), .ZN(n10326)
         );
  nd02d1 U10512 ( .A1(images_bus[364]), .A2(n11752), .ZN(n6313) );
  nd02d1 U10513 ( .A1(images_bus[382]), .A2(images_bus[381]), .ZN(n6594) );
  nd03d1 U10514 ( .A1(n4568), .A2(images_bus[19]), .A3(N8198), .ZN(n10459) );
  nd02d1 U10516 ( .A1(n5414), .A2(images_bus[280]), .ZN(n6612) );
  nd02d1 U10517 ( .A1(images_bus[278]), .A2(n3557), .ZN(n12030) );
  nd02d1 U10518 ( .A1(images_bus[274]), .A2(images_bus[273]), .ZN(n9620) );
  nd03d1 U10519 ( .A1(n11430), .A2(n6139), .A3(images_bus[96]), .ZN(n7572) );
  nd02d1 U10520 ( .A1(n11615), .A2(images_bus[243]), .ZN(n11613) );
  nd02d1 U10521 ( .A1(images_bus[256]), .A2(n3571), .ZN(n11253) );
  nr02d1 U10522 ( .A1(n5455), .A2(n12157), .ZN(n11726) );
  nd02d1 U10523 ( .A1(images_bus[204]), .A2(n9627), .ZN(n9163) );
  nd02d1 U10524 ( .A1(images_bus[366]), .A2(n11753), .ZN(n10931) );
  nd02d1 U10525 ( .A1(images_bus[443]), .A2(n8730), .ZN(n11062) );
  nd03d1 U10526 ( .A1(n4330), .A2(images_bus[55]), .A3(n8221), .ZN(n6725) );
  nd03d1 U10528 ( .A1(n11605), .A2(images_bus[235]), .A3(N11271), .ZN(n6088)
         );
  nd02d1 U10530 ( .A1(images_bus[481]), .A2(images_bus[480]), .ZN(n8830) );
  nd02d1 U10532 ( .A1(n4485), .A2(images_bus[292]), .ZN(n5386) );
  nd03d1 U10533 ( .A1(N13810), .A2(n11989), .A3(images_bus[395]), .ZN(n10984)
         );
  nd03d1 U10534 ( .A1(n5071), .A2(n3873), .A3(images_bus[213]), .ZN(n6960) );
  nd02d1 U10535 ( .A1(images_bus[143]), .A2(n5077), .ZN(n5786) );
  nd02d1 U10536 ( .A1(images_bus[351]), .A2(n6277), .ZN(n8072) );
  nd03d1 U10537 ( .A1(images_bus[254]), .A2(n11622), .A3(images_bus[255]), 
        .ZN(n8463) );
  nd03d1 U10538 ( .A1(n5717), .A2(images_bus[369]), .A3(n5481), .ZN(n5493) );
  nd03d1 U10539 ( .A1(images_bus[336]), .A2(n9347), .A3(n4985), .ZN(n9352) );
  nd03d1 U10540 ( .A1(N11451), .A2(n3793), .A3(images_bus[247]), .ZN(n10746)
         );
  nd03d1 U10543 ( .A1(N14450), .A2(n3115), .A3(images_bus[435]), .ZN(n11838)
         );
  nd03d1 U10544 ( .A1(n4182), .A2(images_bus[73]), .A3(N8896), .ZN(n9012) );
  nd03d1 U10545 ( .A1(n4305), .A2(images_bus[375]), .A3(n9399), .ZN(n9405) );
  nd03d1 U10546 ( .A1(n3876), .A2(images_bus[209]), .A3(N10881), .ZN(n8410) );
  nd03d1 U10548 ( .A1(n3802), .A2(n5939), .A3(images_bus[241]), .ZN(n5321) );
  nd03d1 U10549 ( .A1(n4985), .A2(images_bus[339]), .A3(n5452), .ZN(n5454) );
  nd03d1 U10550 ( .A1(images_bus[119]), .A2(n4322), .A3(n9069), .ZN(n9077) );
  nd03d1 U10552 ( .A1(n9199), .A2(images_bus[229]), .A3(N11181), .ZN(n5289) );
  nd03d1 U10553 ( .A1(images_bus[119]), .A2(n4099), .A3(images_bus[120]), .ZN(
        n6823) );
  inv0d0 U10554 ( .I(n2610), .ZN(N8445) );
  nd02d1 U10555 ( .A1(images_bus[193]), .A2(images_bus[192]), .ZN(n11561) );
  nd03d1 U10556 ( .A1(n4470), .A2(n5192), .A3(images_bus[175]), .ZN(n8091) );
  nd03d1 U10557 ( .A1(n4180), .A2(images_bus[77]), .A3(N8952), .ZN(n6667) );
  nd03d1 U10558 ( .A1(n3277), .A2(n12165), .A3(n6295), .ZN(n6298) );
  nd03d1 U10559 ( .A1(n6271), .A2(images_bus[350]), .A3(images_bus[351]), .ZN(
        n7147) );
  nr02d1 U10560 ( .A1(n9071), .A2(images_bus[117]), .ZN(n9066) );
  nd03d1 U10561 ( .A1(n3122), .A2(n6467), .A3(n3072), .ZN(n6463) );
  inv0d0 U10562 ( .I(n6568), .ZN(n3078) );
  nr02d1 U10563 ( .A1(n7236), .A2(images_bus[399]), .ZN(n4673) );
  nd02d1 U10564 ( .A1(images_bus[429]), .A2(n3122), .ZN(n8704) );
  nd02d1 U10565 ( .A1(images_bus[374]), .A2(images_bus[373]), .ZN(n9606) );
  nd03d1 U10566 ( .A1(n3930), .A2(n10638), .A3(n8356), .ZN(n10636) );
  nd02d1 U10567 ( .A1(images_bus[402]), .A2(images_bus[401]), .ZN(n6402) );
  nd03d1 U10568 ( .A1(n4179), .A2(n7450), .A3(images_bus[81]), .ZN(n6764) );
  inv0d0 U10569 ( .I(n2251), .ZN(n2254) );
  nd02d1 U10570 ( .A1(images_bus[161]), .A2(images_bus[160]), .ZN(n10413) );
  nd03d1 U10571 ( .A1(images_bus[164]), .A2(images_bus[163]), .A3(n4719), .ZN(
        n8093) );
  nr02d1 U10573 ( .A1(n6198), .A2(images_bus[319]), .ZN(n4527) );
  nd02d1 U10574 ( .A1(images_bus[95]), .A2(images_bus[94]), .ZN(n6774) );
  nd03d1 U10576 ( .A1(images_bus[271]), .A2(n3563), .A3(N11826), .ZN(n7762) );
  nd02d1 U10577 ( .A1(images_bus[166]), .A2(images_bus[165]), .ZN(n6885) );
  nd03d1 U10578 ( .A1(N15570), .A2(n11953), .A3(images_bus[505]), .ZN(n11955)
         );
  nd03d1 U10580 ( .A1(images_bus[222]), .A2(n3810), .A3(images_bus[223]), .ZN(
        n11586) );
  nd03d1 U10581 ( .A1(images_bus[17]), .A2(images_bus[16]), .A3(images_bus[18]), .ZN(n7473) );
  nd02d1 U10582 ( .A1(images_bus[461]), .A2(n6279), .ZN(n8767) );
  nd03d1 U10583 ( .A1(images_bus[150]), .A2(n4048), .A3(images_bus[151]), .ZN(
        n5099) );
  nd02d1 U10584 ( .A1(images_bus[449]), .A2(n3010), .ZN(n11852) );
  nd03d1 U10585 ( .A1(images_bus[346]), .A2(n12004), .A3(images_bus[347]), 
        .ZN(n8572) );
  nd02d1 U10586 ( .A1(n9613), .A2(images_bus[322]), .ZN(n8074) );
  nd03d1 U10587 ( .A1(images_bus[274]), .A2(n5362), .A3(images_bus[275]), .ZN(
        n10780) );
  nd03d1 U10588 ( .A1(n4042), .A2(images_bus[154]), .A3(N10056), .ZN(n9847) );
  nd03d1 U10589 ( .A1(n8900), .A2(images_bus[7]), .A3(N8064), .ZN(n8129) );
  nd02d1 U10590 ( .A1(images_bus[426]), .A2(images_bus[425]), .ZN(n8694) );
  nd02d1 U10591 ( .A1(images_bus[230]), .A2(images_bus[229]), .ZN(n9197) );
  nd02d1 U10592 ( .A1(n10069), .A2(images_bus[331]), .ZN(n10063) );
  nd02d1 U10593 ( .A1(images_bus[460]), .A2(images_bus[459]), .ZN(n8759) );
  nd02d1 U10594 ( .A1(images_bus[312]), .A2(images_bus[311]), .ZN(n7395) );
  nd02d1 U10595 ( .A1(n4411), .A2(images_bus[431]), .ZN(n6468) );
  nd02d1 U10596 ( .A1(images_bus[74]), .A2(images_bus[73]), .ZN(n5827) );
  nd02d1 U10597 ( .A1(images_bus[115]), .A2(n6547), .ZN(n8873) );
  nd02d1 U10598 ( .A1(images_bus[65]), .A2(images_bus[64]), .ZN(n5803) );
  nd03d1 U10599 ( .A1(n5729), .A2(images_bus[419]), .A3(n6574), .ZN(n6444) );
  nd02d1 U10600 ( .A1(images_bus[194]), .A2(n6013), .ZN(n9903) );
  nd02d1 U10601 ( .A1(images_bus[219]), .A2(n11583), .ZN(n8424) );
  nd02d1 U10602 ( .A1(images_bus[469]), .A2(n6212), .ZN(n11880) );
  nd03d1 U10604 ( .A1(images_bus[324]), .A2(images_bus[323]), .A3(n6205), .ZN(
        n6208) );
  nd02d1 U10605 ( .A1(n10060), .A2(images_bus[327]), .ZN(n10064) );
  nd02d1 U10606 ( .A1(images_bus[480]), .A2(images_bus[479]), .ZN(n11903) );
  nd02d1 U10607 ( .A1(images_bus[427]), .A2(n6556), .ZN(n7954) );
  nd02d1 U10608 ( .A1(images_bus[227]), .A2(n6621), .ZN(n5754) );
  nd02d1 U10609 ( .A1(images_bus[406]), .A2(n3235), .ZN(n6417) );
  nd02d1 U10610 ( .A1(images_bus[430]), .A2(images_bus[429]), .ZN(n6573) );
  nd02d1 U10611 ( .A1(images_bus[8]), .A2(n5714), .ZN(n8903) );
  nr02d1 U10612 ( .A1(n12127), .A2(n10596), .ZN(n10599) );
  nd02d1 U10613 ( .A1(images_bus[252]), .A2(images_bus[251]), .ZN(n5350) );
  nd02d1 U10614 ( .A1(images_bus[355]), .A2(n6601), .ZN(n4591) );
  nd02d1 U10615 ( .A1(images_bus[330]), .A2(images_bus[329]), .ZN(n5726) );
  nd03d1 U10616 ( .A1(n5406), .A2(images_bus[315]), .A3(n5417), .ZN(n5421) );
  nd02d1 U10617 ( .A1(images_bus[179]), .A2(n6543), .ZN(n7427) );
  nd03d1 U10618 ( .A1(images_bus[486]), .A2(n10292), .A3(images_bus[487]), 
        .ZN(n10298) );
  nd02d1 U10619 ( .A1(images_bus[454]), .A2(n3006), .ZN(n10230) );
  nd02d1 U10620 ( .A1(images_bus[88]), .A2(n11423), .ZN(n7561) );
  nd02d1 U10621 ( .A1(images_bus[276]), .A2(images_bus[275]), .ZN(n5742) );
  nd02d1 U10622 ( .A1(images_bus[11]), .A2(n4832), .ZN(n10430) );
  nd02d1 U10623 ( .A1(images_bus[444]), .A2(images_bus[443]), .ZN(n7974) );
  nd03d1 U10624 ( .A1(n4052), .A2(images_bus[144]), .A3(N9906), .ZN(n10609) );
  nd02d1 U10625 ( .A1(n10332), .A2(images_bus[503]), .ZN(n10334) );
  nd02d1 U10627 ( .A1(n9287), .A2(images_bus[295]), .ZN(n9290) );
  nd02d1 U10628 ( .A1(images_bus[78]), .A2(images_bus[77]), .ZN(n11407) );
  nd02d1 U10629 ( .A1(images_bus[162]), .A2(n3967), .ZN(n6874) );
  nd03d1 U10630 ( .A1(images_bus[41]), .A2(n6702), .A3(n11346), .ZN(n11352) );
  nd02d1 U10631 ( .A1(n5442), .A2(images_bus[152]), .ZN(n7434) );
  nd02d1 U10632 ( .A1(images_bus[438]), .A2(images_bus[437]), .ZN(n5700) );
  nd02d1 U10633 ( .A1(n7135), .A2(n11724), .ZN(n4566) );
  nd02d1 U10634 ( .A1(images_bus[380]), .A2(n9605), .ZN(n9406) );
  nd02d1 U10635 ( .A1(images_bus[129]), .A2(images_bus[128]), .ZN(n5054) );
  nr02d1 U10636 ( .A1(n8621), .A2(images_bus[387]), .ZN(n4642) );
  nd03d1 U10637 ( .A1(n6663), .A2(images_bus[74]), .A3(n4220), .ZN(n8250) );
  inv0d0 U10639 ( .I(n9069), .ZN(n4135) );
  nd02d1 U10640 ( .A1(images_bus[381]), .A2(n10958), .ZN(n7209) );
  nd03d1 U10641 ( .A1(n5061), .A2(images_bus[279]), .A3(n9619), .ZN(n5741) );
  nd03d1 U10642 ( .A1(images_bus[13]), .A2(n4819), .A3(N8129), .ZN(n9664) );
  nd03d1 U10643 ( .A1(n9697), .A2(n8119), .A3(images_bus[37]), .ZN(n10486) );
  nd02d1 U10645 ( .A1(images_bus[448]), .A2(n8738), .ZN(n11849) );
  nd03d1 U10646 ( .A1(N14962), .A2(n11970), .A3(images_bus[467]), .ZN(n11877)
         );
  nd02d1 U10647 ( .A1(n10321), .A2(images_bus[499]), .ZN(n10328) );
  nd02d1 U10648 ( .A1(images_bus[6]), .A2(n4858), .ZN(n9657) );
  nd03d1 U10649 ( .A1(images_bus[129]), .A2(n11473), .A3(images_bus[130]), 
        .ZN(n5961) );
  nr02d1 U10650 ( .A1(n9235), .A2(images_bus[253]), .ZN(n7020) );
  nr02d1 U10651 ( .A1(n7857), .A2(images_bus[359]), .ZN(n4598) );
  nd03d1 U10652 ( .A1(n3475), .A2(n6922), .A3(images_bus[291]), .ZN(n6172) );
  nd03d1 U10654 ( .A1(images_bus[140]), .A2(images_bus[139]), .A3(n11491), 
        .ZN(n11496) );
  nd03d1 U10655 ( .A1(N13890), .A2(n3200), .A3(images_bus[400]), .ZN(n11984)
         );
  nd03d1 U10656 ( .A1(images_bus[408]), .A2(n8658), .A3(images_bus[409]), .ZN(
        n7368) );
  nr02d1 U10657 ( .A1(n6372), .A2(images_bus[389]), .ZN(n4652) );
  nd03d1 U10658 ( .A1(images_bus[438]), .A2(n10201), .A3(images_bus[439]), 
        .ZN(n10210) );
  nd03d1 U10659 ( .A1(n4315), .A2(images_bus[215]), .A3(n9176), .ZN(n9178) );
  nd02d1 U10660 ( .A1(images_bus[163]), .A2(n3966), .ZN(n10632) );
  nr02d1 U10661 ( .A1(n5715), .A2(n12125), .ZN(n7345) );
  nd03d1 U10662 ( .A1(images_bus[6]), .A2(n8897), .A3(images_bus[7]), .ZN(
        n8901) );
  nd03d1 U10663 ( .A1(n11338), .A2(images_bus[32]), .A3(N8354), .ZN(n10478) );
  nd03d1 U10664 ( .A1(images_bus[198]), .A2(n9901), .A3(images_bus[199]), .ZN(
        n9904) );
  nr02d1 U10666 ( .A1(n6987), .A2(images_bus[235]), .ZN(n9949) );
  nd03d1 U10667 ( .A1(n9081), .A2(n4966), .A3(images_bus[125]), .ZN(n9811) );
  nd03d1 U10668 ( .A1(images_bus[214]), .A2(n3870), .A3(N10956), .ZN(n5248) );
  nd02d1 U10670 ( .A1(images_bus[324]), .A2(n11696), .ZN(n10861) );
  nd02d1 U10673 ( .A1(n9913), .A2(images_bus[207]), .ZN(n9914) );
  nd03d1 U10674 ( .A1(n4309), .A2(images_bus[274]), .A3(n3519), .ZN(n6150) );
  nd03d1 U10675 ( .A1(n3965), .A2(images_bus[164]), .A3(N10206), .ZN(n10630)
         );
  nd03d1 U10676 ( .A1(n4656), .A2(images_bus[359]), .A3(n9381), .ZN(n9385) );
  nd02d1 U10677 ( .A1(images_bus[389]), .A2(n3244), .ZN(n9422) );
  nd02d1 U10678 ( .A1(images_bus[224]), .A2(images_bus[223]), .ZN(n6622) );
  nd02d1 U10679 ( .A1(images_bus[362]), .A2(n7384), .ZN(n5485) );
  nd02d1 U10680 ( .A1(images_bus[385]), .A2(images_bus[384]), .ZN(n6367) );
  nr02d1 U10681 ( .A1(n6777), .A2(n10411), .ZN(n9880) );
  nd03d1 U10682 ( .A1(images_bus[416]), .A2(n8681), .A3(images_bus[417]), .ZN(
        n8673) );
  nd03d1 U10683 ( .A1(images_bus[159]), .A2(n7648), .A3(N10131), .ZN(n5981) );
  nd03d1 U10684 ( .A1(images_bus[57]), .A2(n12071), .A3(N8679), .ZN(n8979) );
  nd02d1 U10685 ( .A1(images_bus[440]), .A2(n11055), .ZN(n11058) );
  nd03d1 U10686 ( .A1(n10426), .A2(images_bus[42]), .A3(N8484), .ZN(n7502) );
  nd02d1 U10687 ( .A1(n7536), .A2(images_bus[75]), .ZN(n8111) );
  nd02d1 U10688 ( .A1(images_bus[418]), .A2(n8680), .ZN(n11980) );
  nd03d1 U10689 ( .A1(n9023), .A2(n6661), .A3(n9025), .ZN(n9024) );
  inv0d0 U10691 ( .I(n9031), .ZN(n4141) );
  nd03d1 U10692 ( .A1(n4179), .A2(images_bus[79]), .A3(N8980), .ZN(n10537) );
  nd02d1 U10693 ( .A1(n9321), .A2(images_bus[319]), .ZN(n9612) );
  nd02d1 U10694 ( .A1(n5252), .A2(images_bus[357]), .ZN(n6294) );
  nd02d1 U10695 ( .A1(n3191), .A2(n12171), .ZN(n8635) );
  nd03d1 U10696 ( .A1(N11714), .A2(n3534), .A3(images_bus[264]), .ZN(n8473) );
  nd03d1 U10697 ( .A1(images_bus[494]), .A2(n10310), .A3(images_bus[495]), 
        .ZN(n10347) );
  nd02d1 U10698 ( .A1(images_bus[265]), .A2(images_bus[264]), .ZN(n9982) );
  nd03d1 U10699 ( .A1(images_bus[111]), .A2(n12064), .A3(N9428), .ZN(n7585) );
  nd03d1 U10701 ( .A1(n3802), .A2(images_bus[239]), .A3(N11331), .ZN(n9953) );
  nd02d1 U10702 ( .A1(n9272), .A2(images_bus[287]), .ZN(n9616) );
  nr02d1 U10704 ( .A1(n6330), .A2(n10415), .ZN(n9832) );
  nd03d1 U10705 ( .A1(n3350), .A2(n4537), .A3(images_bus[324]), .ZN(n4541) );
  nd03d1 U10706 ( .A1(images_bus[367]), .A2(n3289), .A3(N13362), .ZN(n10932)
         );
  nd03d1 U10707 ( .A1(n2868), .A2(n12166), .A3(n11190), .ZN(n8803) );
  nr02d1 U10708 ( .A1(n10097), .A2(images_bus[367]), .ZN(n6317) );
  nd02d1 U10710 ( .A1(images_bus[402]), .A2(n11983), .ZN(n9436) );
  nd02d1 U10712 ( .A1(images_bus[401]), .A2(images_bus[400]), .ZN(n10389) );
  nr02d1 U10714 ( .A1(n6240), .A2(n10394), .ZN(n10035) );
  nd02d1 U10715 ( .A1(images_bus[438]), .A2(n11978), .ZN(n11973) );
  nd03d1 U10716 ( .A1(images_bus[268]), .A2(images_bus[267]), .A3(n5647), .ZN(
        n8482) );
  nd02d1 U10717 ( .A1(images_bus[449]), .A2(images_bus[448]), .ZN(n10371) );
  nd03d1 U10718 ( .A1(n5997), .A2(images_bus[358]), .A3(n7853), .ZN(n7855) );
  nd03d1 U10719 ( .A1(images_bus[169]), .A2(n9862), .A3(images_bus[168]), .ZN(
        n9873) );
  nd02d1 U10720 ( .A1(n9748), .A2(images_bus[71]), .ZN(n9744) );
  nd03d1 U10724 ( .A1(images_bus[57]), .A2(images_bus[56]), .A3(images_bus[58]), .ZN(n8977) );
  nd03d1 U10725 ( .A1(n4500), .A2(images_bus[303]), .A3(n4994), .ZN(n4519) );
  nd02d1 U10726 ( .A1(images_bus[422]), .A2(n9459), .ZN(n11022) );
  nd02d1 U10729 ( .A1(images_bus[466]), .A2(images_bus[465]), .ZN(n11878) );
  nd02d1 U10730 ( .A1(images_bus[239]), .A2(n4457), .ZN(n8078) );
  nd03d1 U10731 ( .A1(images_bus[406]), .A2(n10149), .A3(images_bus[407]), 
        .ZN(n10151) );
  nd02d1 U10732 ( .A1(images_bus[384]), .A2(n10961), .ZN(n10965) );
  nd03d1 U10734 ( .A1(images_bus[152]), .A2(n4037), .A3(N10026), .ZN(n5102) );
  nd03d1 U10735 ( .A1(images_bus[126]), .A2(n4057), .A3(N9638), .ZN(n10587) );
  nd03d1 U10736 ( .A1(n4437), .A2(images_bus[304]), .A3(n3489), .ZN(n7080) );
  nd03d1 U10737 ( .A1(n3879), .A2(images_bus[199]), .A3(N10731), .ZN(n11571)
         );
  nd02d1 U10738 ( .A1(images_bus[233]), .A2(n7153), .ZN(n9625) );
  nd03d1 U10739 ( .A1(images_bus[102]), .A2(n10420), .A3(images_bus[103]), 
        .ZN(n9786) );
  nd03d1 U10740 ( .A1(images_bus[7]), .A2(n4847), .A3(images_bus[8]), .ZN(
        n11311) );
  nd03d1 U10741 ( .A1(n4201), .A2(images_bus[64]), .A3(N8770), .ZN(n11390) );
  nd03d1 U10742 ( .A1(images_bus[220]), .A2(n3864), .A3(images_bus[221]), .ZN(
        n6966) );
  nr02d1 U10743 ( .A1(n6310), .A2(n10408), .ZN(n9950) );
  nd03d1 U10744 ( .A1(n4604), .A2(images_bus[15]), .A3(N8151), .ZN(n10453) );
  nd03d1 U10745 ( .A1(n5734), .A2(images_bus[323]), .A3(n3338), .ZN(n5439) );
  nd02d1 U10746 ( .A1(images_bus[20]), .A2(images_bus[19]), .ZN(n8888) );
  nd03d1 U10748 ( .A1(N13602), .A2(n3169), .A3(images_bus[382]), .ZN(n11225)
         );
  nd02d1 U10749 ( .A1(images_bus[164]), .A2(n9634), .ZN(n9123) );
  nd02d1 U10750 ( .A1(images_bus[108]), .A2(n9641), .ZN(n9054) );
  nd03d1 U10751 ( .A1(N14770), .A2(n2951), .A3(images_bus[455]), .ZN(n11860)
         );
  nd02d1 U10752 ( .A1(n6496), .A2(n9642), .ZN(n9031) );
  nd03d1 U10753 ( .A1(n4994), .A2(images_bus[303]), .A3(n11669), .ZN(n11685)
         );
  nd02d1 U10754 ( .A1(images_bus[306]), .A2(images_bus[305]), .ZN(n7087) );
  nd02d1 U10755 ( .A1(n10157), .A2(images_bus[411]), .ZN(n10387) );
  nd03d1 U10756 ( .A1(images_bus[224]), .A2(n3736), .A3(N11106), .ZN(n5280) );
  nd02d1 U10758 ( .A1(images_bus[104]), .A2(n8879), .ZN(n8878) );
  nd03d1 U10760 ( .A1(images_bus[2]), .A2(images_bus[1]), .A3(N8016), .ZN(
        n6680) );
  nd03d1 U10762 ( .A1(images_bus[17]), .A2(n4590), .A3(N8174), .ZN(n9671) );
  nd02d1 U10763 ( .A1(n6661), .A2(images_bus[87]), .ZN(n8109) );
  nd03d1 U10764 ( .A1(images_bus[220]), .A2(n3864), .A3(N11046), .ZN(n5264) );
  nd02d1 U10765 ( .A1(images_bus[332]), .A2(n9611), .ZN(n9338) );
  nd03d1 U10766 ( .A1(images_bus[424]), .A2(n9471), .A3(images_bus[425]), .ZN(
        n9469) );
  nd02d1 U10768 ( .A1(images_bus[490]), .A2(n10300), .ZN(n10351) );
  nd03d1 U10769 ( .A1(n11333), .A2(images_bus[25]), .A3(N8270), .ZN(n8165) );
  inv0d0 U10770 ( .I(n2642), .ZN(N8270) );
  inv0d0 U10771 ( .I(n2641), .ZN(n2643) );
  nd02d1 U10774 ( .A1(images_bus[38]), .A2(n4276), .ZN(n6696) );
  nd02d1 U10775 ( .A1(images_bus[133]), .A2(images_bus[132]), .ZN(n10416) );
  nd02d1 U10776 ( .A1(images_bus[26]), .A2(n10427), .ZN(n9681) );
  nd02d1 U10777 ( .A1(n3995), .A2(images_bus[127]), .ZN(n9640) );
  nd02d1 U10778 ( .A1(n6795), .A2(n10418), .ZN(n9801) );
  nd02d1 U10779 ( .A1(n9337), .A2(images_bus[327]), .ZN(n9341) );
  nd02d1 U10780 ( .A1(images_bus[502]), .A2(n4297), .ZN(n9579) );
  nd02d1 U10781 ( .A1(images_bus[434]), .A2(n3116), .ZN(n9477) );
  nd02d1 U10782 ( .A1(images_bus[271]), .A2(n9246), .ZN(n7406) );
  nd02d1 U10783 ( .A1(images_bus[277]), .A2(images_bus[276]), .ZN(n10397) );
  nd02d1 U10784 ( .A1(images_bus[499]), .A2(n11937), .ZN(n11159) );
  nd02d1 U10785 ( .A1(images_bus[299]), .A2(n5642), .ZN(n8512) );
  nd02d1 U10786 ( .A1(images_bus[72]), .A2(images_bus[73]), .ZN(n9011) );
  nd02d1 U10787 ( .A1(images_bus[165]), .A2(images_bus[164]), .ZN(n10412) );
  nd03d1 U10788 ( .A1(images_bus[167]), .A2(images_bus[166]), .A3(n8350), .ZN(
        n8355) );
  nd02d1 U10789 ( .A1(images_bus[147]), .A2(n6544), .ZN(n8097) );
  nd02d1 U10790 ( .A1(images_bus[445]), .A2(n6157), .ZN(n9496) );
  nd03d1 U10791 ( .A1(images_bus[230]), .A2(n9946), .A3(images_bus[231]), .ZN(
        n9941) );
  nd02d1 U10792 ( .A1(images_bus[161]), .A2(n9857), .ZN(n5121) );
  nd02d1 U10793 ( .A1(images_bus[464]), .A2(n11200), .ZN(n11099) );
  nd03d1 U10794 ( .A1(n5061), .A2(images_bus[277]), .A3(n8487), .ZN(n8489) );
  nd03d1 U10795 ( .A1(n10194), .A2(n6556), .A3(images_bus[429]), .ZN(n10193)
         );
  nd02d1 U10796 ( .A1(images_bus[286]), .A2(images_bus[285]), .ZN(n6611) );
  nd02d1 U10797 ( .A1(images_bus[54]), .A2(n4331), .ZN(n11371) );
  nd02d1 U10798 ( .A1(images_bus[266]), .A2(images_bus[265]), .ZN(n8475) );
  nd02d1 U10799 ( .A1(images_bus[358]), .A2(images_bus[357]), .ZN(n7158) );
  nd03d1 U10800 ( .A1(images_bus[359]), .A2(images_bus[358]), .A3(n8591), .ZN(
        n8592) );
  nd02d1 U10801 ( .A1(images_bus[302]), .A2(images_bus[301]), .ZN(n9299) );
  nd02d1 U10802 ( .A1(images_bus[98]), .A2(n5888), .ZN(n11434) );
  nd02d1 U10803 ( .A1(images_bus[178]), .A2(images_bus[177]), .ZN(n8370) );
  nd02d1 U10804 ( .A1(images_bus[300]), .A2(n3462), .ZN(n10023) );
  nd02d1 U10805 ( .A1(images_bus[231]), .A2(n3808), .ZN(n5292) );
  nd02d1 U10806 ( .A1(images_bus[69]), .A2(n11392), .ZN(n9000) );
  nd03d1 U10807 ( .A1(images_bus[208]), .A2(n9914), .A3(images_bus[209]), .ZN(
        n9915) );
  nd03d1 U10808 ( .A1(images_bus[58]), .A2(n9729), .A3(images_bus[59]), .ZN(
        n9732) );
  nd02d1 U10809 ( .A1(images_bus[477]), .A2(n6155), .ZN(n7998) );
  nd02d1 U10810 ( .A1(images_bus[282]), .A2(images_bus[281]), .ZN(n12033) );
  nd02d1 U10811 ( .A1(images_bus[143]), .A2(n4054), .ZN(n11503) );
  nd02d1 U10812 ( .A1(images_bus[131]), .A2(n4056), .ZN(n5048) );
  nd02d1 U10813 ( .A1(images_bus[149]), .A2(n4050), .ZN(n6858) );
  nd03d1 U10815 ( .A1(n5910), .A2(images_bus[401]), .A3(n7229), .ZN(n7231) );
  nd02d1 U10816 ( .A1(images_bus[417]), .A2(n10386), .ZN(n7923) );
  nd02d1 U10818 ( .A1(images_bus[21]), .A2(n11324), .ZN(n8159) );
  nd02d1 U10819 ( .A1(n4742), .A2(images_bus[131]), .ZN(n8100) );
  nd02d1 U10820 ( .A1(images_bus[99]), .A2(images_bus[100]), .ZN(n11440) );
  nd02d1 U10821 ( .A1(images_bus[132]), .A2(n9638), .ZN(n6848) );
  nd02d1 U10822 ( .A1(images_bus[144]), .A2(n5082), .ZN(n9636) );
  nd02d1 U10823 ( .A1(images_bus[54]), .A2(n10503), .ZN(n10507) );
  nd02d1 U10824 ( .A1(images_bus[70]), .A2(images_bus[69]), .ZN(n5815) );
  nd03d1 U10825 ( .A1(n7422), .A2(images_bus[196]), .A3(n3886), .ZN(n11565) );
  nr02d1 U10826 ( .A1(n6291), .A2(n12171), .ZN(n4964) );
  nd02d1 U10827 ( .A1(n10185), .A2(images_bus[427]), .ZN(n10194) );
  nd02d1 U10828 ( .A1(n9840), .A2(images_bus[151]), .ZN(n9845) );
  nd02d1 U10829 ( .A1(images_bus[26]), .A2(n10464), .ZN(n10467) );
  nd03d1 U10830 ( .A1(N11602), .A2(n3527), .A3(images_bus[257]), .ZN(n11252)
         );
  nd03d1 U10831 ( .A1(n4168), .A2(n4169), .A3(n9771), .ZN(n9768) );
  nd02d1 U10834 ( .A1(images_bus[16]), .A2(n10447), .ZN(n10449) );
  nd03d1 U10835 ( .A1(images_bus[207]), .A2(images_bus[204]), .A3(n4462), .ZN(
        n7419) );
  nd02d1 U10836 ( .A1(images_bus[264]), .A2(n10765), .ZN(n10768) );
  nd02d1 U10837 ( .A1(images_bus[416]), .A2(n7367), .ZN(n7266) );
  nd02d1 U10839 ( .A1(n8440), .A2(images_bus[237]), .ZN(n6988) );
  nd02d1 U10840 ( .A1(images_bus[234]), .A2(n10718), .ZN(n10720) );
  nd03d1 U10841 ( .A1(images_bus[312]), .A2(n9311), .A3(n5406), .ZN(n9314) );
  nd03d1 U10842 ( .A1(n4510), .A2(images_bus[76]), .A3(n4209), .ZN(n7545) );
  nd02d1 U10843 ( .A1(images_bus[254]), .A2(n10748), .ZN(n10752) );
  nd03d1 U10844 ( .A1(n2917), .A2(n6279), .A3(images_bus[463]), .ZN(n10364) );
  nd02d1 U10845 ( .A1(n7914), .A2(images_bus[415]), .ZN(n7920) );
  nd03d1 U10846 ( .A1(images_bus[184]), .A2(n9143), .A3(n5435), .ZN(n9149) );
  nd02d1 U10847 ( .A1(images_bus[430]), .A2(n11040), .ZN(n11213) );
  nd03d1 U10848 ( .A1(images_bus[152]), .A2(n9845), .A3(images_bus[153]), .ZN(
        n9842) );
  nd03d1 U10849 ( .A1(n10328), .A2(n4297), .A3(images_bus[500]), .ZN(n10323)
         );
  nd02d1 U10852 ( .A1(images_bus[98]), .A2(n9785), .ZN(n9782) );
  nd02d1 U10854 ( .A1(images_bus[86]), .A2(n10422), .ZN(n9763) );
  nd03d1 U10855 ( .A1(n4444), .A2(images_bus[264]), .A3(n3510), .ZN(n11642) );
  nd03d1 U10856 ( .A1(n4444), .A2(images_bus[264]), .A3(n4681), .ZN(n4452) );
  nd03d1 U10857 ( .A1(images_bus[170]), .A2(n9873), .A3(images_bus[171]), .ZN(
        n9868) );
  nd03d1 U10858 ( .A1(n10837), .A2(n10838), .A3(n3454), .ZN(n10836) );
  nd02d1 U10859 ( .A1(images_bus[41]), .A2(n11294), .ZN(n10488) );
  nd02d1 U10860 ( .A1(images_bus[490]), .A2(n5604), .ZN(n8829) );
  nd02d1 U10861 ( .A1(n5714), .A2(n11299), .ZN(n10440) );
  nd02d1 U10862 ( .A1(n6793), .A2(images_bus[104]), .ZN(n6796) );
  nd03d1 U10863 ( .A1(n4323), .A2(images_bus[88]), .A3(n11419), .ZN(n11422) );
  nd02d1 U10864 ( .A1(n9891), .A2(images_bus[191]), .ZN(n9894) );
  nd02d1 U10865 ( .A1(images_bus[430]), .A2(n10193), .ZN(n10187) );
  nd02d1 U10868 ( .A1(n10123), .A2(images_bus[391]), .ZN(n10127) );
  nd02d1 U10869 ( .A1(images_bus[257]), .A2(images_bus[256]), .ZN(n10405) );
  nd03d1 U10870 ( .A1(images_bus[196]), .A2(images_bus[195]), .A3(n5199), .ZN(
        n5764) );
  nd02d1 U10871 ( .A1(images_bus[110]), .A2(n10419), .ZN(n9797) );
  nd02d1 U10872 ( .A1(images_bus[149]), .A2(n11272), .ZN(n10611) );
  nd02d1 U10873 ( .A1(images_bus[210]), .A2(n9915), .ZN(n9918) );
  nd02d1 U10874 ( .A1(n9743), .A2(images_bus[67]), .ZN(n9745) );
  nd02d1 U10875 ( .A1(images_bus[184]), .A2(n10650), .ZN(n10653) );
  inv0d0 U10876 ( .I(n11264), .ZN(n3906) );
  nd02d1 U10877 ( .A1(n3482), .A2(images_bus[315]), .ZN(n10040) );
  nd02d1 U10879 ( .A1(n6543), .A2(n9630), .ZN(n9137) );
  nd02d1 U10880 ( .A1(images_bus[364]), .A2(n9608), .ZN(n9391) );
  nd02d1 U10882 ( .A1(images_bus[396]), .A2(n4416), .ZN(n10135) );
  nd02d1 U10883 ( .A1(images_bus[184]), .A2(images_bus[185]), .ZN(n9886) );
  nd02d1 U10884 ( .A1(images_bus[66]), .A2(n11288), .ZN(n10521) );
  nd02d1 U10885 ( .A1(images_bus[379]), .A2(n6664), .ZN(n10112) );
  nd02d1 U10886 ( .A1(images_bus[465]), .A2(n11099), .ZN(n11100) );
  nd02d1 U10887 ( .A1(images_bus[416]), .A2(n7920), .ZN(n7924) );
  nd02d1 U10888 ( .A1(images_bus[360]), .A2(n8592), .ZN(n8589) );
  inv0d0 U10889 ( .I(n11809), .ZN(n3210) );
  inv0d0 U10890 ( .I(n11636), .ZN(n3568) );
  inv0d0 U10891 ( .I(n6255), .ZN(n2801) );
  nd02d1 U10892 ( .A1(images_bus[492]), .A2(n9562), .ZN(n10353) );
  aoim22d1 U10893 ( .A1(n9392), .A2(n3286), .B1(n9393), .B2(n9394), .Z(n9386)
         );
  nd02d1 U10896 ( .A1(n5274), .A2(images_bus[229]), .ZN(n7716) );
  buffd1 U10898 ( .I(num_images[2]), .Z(n1039) );
  buffd1 U10899 ( .I(num_images[2]), .Z(n1040) );
  buffd1 U10900 ( .I(num_images[2]), .Z(n1038) );
  buffd1 U10901 ( .I(num_images[2]), .Z(n1037) );
  buffd1 U10902 ( .I(n1041), .Z(n1086) );
  buffd1 U10903 ( .I(num_images[2]), .Z(n1041) );
  aoim22d1 U10904 ( .A1(n6925), .A2(n6926), .B1(n6927), .B2(n6928), .Z(n6924)
         );
  inv0d0 U10906 ( .I(num_images[6]), .ZN(n1222) );
  inv0d0 U10907 ( .I(num_images[7]), .ZN(n1271) );
  inv0d0 U10908 ( .I(N6867), .ZN(n958) );
  inv0d0 U10909 ( .I(num_images[3]), .ZN(n1088) );
  inv0d0 U10910 ( .I(num_images[4]), .ZN(n1133) );
  inv0d0 U10911 ( .I(num_images[5]), .ZN(n1176) );
  inv0d0 U10912 ( .I(N11556), .ZN(n1372) );
  nr02d0 U10992 ( .A1(n501), .A2(n500), .ZN(n29) );
  an02d0 U10993 ( .A1(n29), .A2(n513), .Z(n392) );
  nr02d0 U10994 ( .A1(n501), .A2(n499), .ZN(n30) );
  an02d0 U10995 ( .A1(n513), .A2(n30), .Z(n391) );
  aoi22d1 U10996 ( .A1(images_bus[229]), .A2(n436), .B1(images_bus[231]), .B2(
        n426), .ZN(n36) );
  nr02d0 U10997 ( .A1(N3973), .A2(N3974), .ZN(n31) );
  an02d0 U10998 ( .A1(n31), .A2(n513), .Z(n394) );
  nr02d0 U10999 ( .A1(n499), .A2(N3974), .ZN(n32) );
  an02d0 U11000 ( .A1(n32), .A2(n513), .Z(n393) );
  aoi22d1 U11001 ( .A1(images_bus[225]), .A2(n455), .B1(images_bus[227]), .B2(
        n445), .ZN(n35) );
  an02d0 U11002 ( .A1(n29), .A2(n512), .Z(n396) );
  an02d0 U11003 ( .A1(n30), .A2(n512), .Z(n395) );
  aoi22d1 U11004 ( .A1(n6621), .A2(n474), .B1(images_bus[230]), .B2(n464), 
        .ZN(n34) );
  an02d0 U11005 ( .A1(n32), .A2(n512), .Z(n397) );
  aoi22d1 U11006 ( .A1(images_bus[224]), .A2(n492), .B1(n6931), .B2(n481), 
        .ZN(n33) );
  nd04d0 U11007 ( .A1(n36), .A2(n35), .A3(n34), .A4(n33), .ZN(n42) );
  aoi22d1 U11008 ( .A1(images_bus[245]), .A2(n436), .B1(images_bus[247]), .B2(
        n426), .ZN(n40) );
  aoi22d1 U11009 ( .A1(images_bus[241]), .A2(n455), .B1(images_bus[243]), .B2(
        n445), .ZN(n39) );
  aoi22d1 U11010 ( .A1(images_bus[244]), .A2(n474), .B1(images_bus[246]), .B2(
        n464), .ZN(n38) );
  aoi22d1 U11011 ( .A1(images_bus[240]), .A2(n492), .B1(images_bus[242]), .B2(
        n481), .ZN(n37) );
  nd04d0 U11012 ( .A1(n40), .A2(n39), .A3(n38), .A4(n37), .ZN(n41) );
  aoi22d1 U11013 ( .A1(n42), .A2(n385), .B1(n41), .B2(n383), .ZN(n77) );
  aoi22d1 U11014 ( .A1(n4698), .A2(n436), .B1(images_bus[199]), .B2(n426), 
        .ZN(n46) );
  aoi22d1 U11015 ( .A1(images_bus[193]), .A2(n455), .B1(images_bus[195]), .B2(
        n445), .ZN(n45) );
  aoi22d1 U11016 ( .A1(images_bus[196]), .A2(n474), .B1(images_bus[198]), .B2(
        n464), .ZN(n44) );
  aoi22d1 U11017 ( .A1(images_bus[192]), .A2(n492), .B1(images_bus[194]), .B2(
        n477), .ZN(n43) );
  nd04d0 U11018 ( .A1(n46), .A2(n45), .A3(n44), .A4(n43), .ZN(n52) );
  aoi22d1 U11019 ( .A1(images_bus[213]), .A2(n436), .B1(images_bus[215]), .B2(
        n426), .ZN(n50) );
  aoi22d1 U11020 ( .A1(images_bus[209]), .A2(n455), .B1(images_bus[211]), .B2(
        n445), .ZN(n49) );
  aoi22d1 U11021 ( .A1(images_bus[212]), .A2(n474), .B1(images_bus[214]), .B2(
        n464), .ZN(n48) );
  aoi22d1 U11022 ( .A1(images_bus[208]), .A2(n492), .B1(images_bus[210]), .B2(
        n479), .ZN(n47) );
  nd04d0 U11023 ( .A1(n50), .A2(n49), .A3(n48), .A4(n47), .ZN(n51) );
  aoi22d1 U11024 ( .A1(n52), .A2(n404), .B1(n51), .B2(n402), .ZN(n76) );
  aoi22d1 U11025 ( .A1(images_bus[237]), .A2(n436), .B1(images_bus[239]), .B2(
        n426), .ZN(n56) );
  aoi22d1 U11026 ( .A1(images_bus[233]), .A2(n455), .B1(images_bus[235]), .B2(
        n445), .ZN(n55) );
  aoi22d1 U11027 ( .A1(images_bus[236]), .A2(n474), .B1(images_bus[238]), .B2(
        n464), .ZN(n54) );
  aoi22d1 U11028 ( .A1(n7153), .A2(n492), .B1(images_bus[234]), .B2(n477), 
        .ZN(n53) );
  nd04d0 U11029 ( .A1(n56), .A2(n55), .A3(n54), .A4(n53), .ZN(n62) );
  aoi22d1 U11030 ( .A1(images_bus[253]), .A2(n436), .B1(images_bus[255]), .B2(
        n426), .ZN(n60) );
  aoi22d1 U11031 ( .A1(images_bus[249]), .A2(n455), .B1(images_bus[251]), .B2(
        n445), .ZN(n59) );
  aoi22d1 U11032 ( .A1(images_bus[252]), .A2(n474), .B1(images_bus[254]), .B2(
        n464), .ZN(n58) );
  aoi22d1 U11033 ( .A1(images_bus[248]), .A2(n492), .B1(images_bus[250]), .B2(
        n477), .ZN(n57) );
  nd04d0 U11034 ( .A1(n60), .A2(n59), .A3(n58), .A4(n57), .ZN(n61) );
  aoi22d1 U11035 ( .A1(n62), .A2(n385), .B1(n61), .B2(n383), .ZN(n74) );
  aoi22d1 U11036 ( .A1(images_bus[205]), .A2(n436), .B1(images_bus[207]), .B2(
        n426), .ZN(n66) );
  aoi22d1 U11037 ( .A1(images_bus[201]), .A2(n455), .B1(images_bus[203]), .B2(
        n445), .ZN(n65) );
  aoi22d1 U11038 ( .A1(images_bus[204]), .A2(n474), .B1(n6324), .B2(n464), 
        .ZN(n64) );
  aoi22d1 U11039 ( .A1(images_bus[200]), .A2(n492), .B1(n6861), .B2(n477), 
        .ZN(n63) );
  nd04d0 U11040 ( .A1(n66), .A2(n65), .A3(n64), .A4(n63), .ZN(n72) );
  aoi22d1 U11041 ( .A1(images_bus[221]), .A2(n436), .B1(images_bus[223]), .B2(
        n426), .ZN(n70) );
  aoi22d1 U11042 ( .A1(images_bus[217]), .A2(n455), .B1(images_bus[219]), .B2(
        n445), .ZN(n69) );
  aoi22d1 U11043 ( .A1(images_bus[220]), .A2(n474), .B1(images_bus[222]), .B2(
        n464), .ZN(n68) );
  aoi22d1 U11044 ( .A1(images_bus[216]), .A2(n492), .B1(n6682), .B2(n477), 
        .ZN(n67) );
  nd04d0 U11045 ( .A1(n70), .A2(n69), .A3(n68), .A4(n67), .ZN(n71) );
  aoi22d1 U11046 ( .A1(n72), .A2(n404), .B1(n71), .B2(n402), .ZN(n73) );
  oaim21d1 U11047 ( .B1(n74), .B2(n73), .A(n955), .ZN(n75) );
  aon211d1 U11048 ( .C1(n77), .C2(n76), .B(n955), .A(n75), .ZN(n124) );
  aoi22d1 U11049 ( .A1(images_bus[165]), .A2(n436), .B1(images_bus[167]), .B2(
        n426), .ZN(n81) );
  aoi22d1 U11050 ( .A1(images_bus[161]), .A2(n455), .B1(images_bus[163]), .B2(
        n445), .ZN(n80) );
  aoi22d1 U11051 ( .A1(images_bus[164]), .A2(n474), .B1(images_bus[166]), .B2(
        n464), .ZN(n79) );
  aoi22d1 U11052 ( .A1(images_bus[160]), .A2(n492), .B1(images_bus[162]), .B2(
        n477), .ZN(n78) );
  nd04d0 U11053 ( .A1(n81), .A2(n80), .A3(n79), .A4(n78), .ZN(n87) );
  aoi22d1 U11054 ( .A1(images_bus[181]), .A2(n435), .B1(images_bus[183]), .B2(
        n425), .ZN(n85) );
  aoi22d1 U11055 ( .A1(images_bus[177]), .A2(n454), .B1(images_bus[179]), .B2(
        n444), .ZN(n84) );
  aoi22d1 U11056 ( .A1(n6543), .A2(n473), .B1(images_bus[182]), .B2(n463), 
        .ZN(n83) );
  aoi22d1 U11057 ( .A1(images_bus[176]), .A2(n491), .B1(images_bus[178]), .B2(
        n477), .ZN(n82) );
  nd04d0 U11058 ( .A1(n85), .A2(n84), .A3(n83), .A4(n82), .ZN(n86) );
  aoi22d1 U11059 ( .A1(n87), .A2(n385), .B1(n86), .B2(n383), .ZN(n122) );
  aoi22d1 U11060 ( .A1(images_bus[133]), .A2(n435), .B1(images_bus[135]), .B2(
        n425), .ZN(n91) );
  aoi22d1 U11061 ( .A1(images_bus[129]), .A2(n454), .B1(images_bus[131]), .B2(
        n444), .ZN(n90) );
  aoi22d1 U11062 ( .A1(images_bus[132]), .A2(n473), .B1(images_bus[134]), .B2(
        n463), .ZN(n89) );
  aoi22d1 U11063 ( .A1(images_bus[128]), .A2(n491), .B1(images_bus[130]), .B2(
        n477), .ZN(n88) );
  nd04d0 U11064 ( .A1(n91), .A2(n90), .A3(n89), .A4(n88), .ZN(n97) );
  aoi22d1 U11065 ( .A1(images_bus[149]), .A2(n435), .B1(images_bus[151]), .B2(
        n425), .ZN(n95) );
  aoi22d1 U11066 ( .A1(images_bus[145]), .A2(n454), .B1(images_bus[147]), .B2(
        n444), .ZN(n94) );
  aoi22d1 U11067 ( .A1(n6544), .A2(n473), .B1(images_bus[150]), .B2(n463), 
        .ZN(n93) );
  aoi22d1 U11068 ( .A1(images_bus[144]), .A2(n491), .B1(images_bus[146]), .B2(
        n478), .ZN(n92) );
  nd04d0 U11069 ( .A1(n95), .A2(n94), .A3(n93), .A4(n92), .ZN(n96) );
  aoi22d1 U11070 ( .A1(n97), .A2(n404), .B1(n96), .B2(n402), .ZN(n121) );
  aoi22d1 U11071 ( .A1(images_bus[173]), .A2(n435), .B1(images_bus[175]), .B2(
        n425), .ZN(n101) );
  aoi22d1 U11072 ( .A1(images_bus[169]), .A2(n454), .B1(images_bus[171]), .B2(
        n444), .ZN(n100) );
  aoi22d1 U11073 ( .A1(images_bus[172]), .A2(n473), .B1(n6328), .B2(n463), 
        .ZN(n99) );
  aoi22d1 U11074 ( .A1(images_bus[168]), .A2(n491), .B1(images_bus[170]), .B2(
        n481), .ZN(n98) );
  nd04d0 U11075 ( .A1(n101), .A2(n100), .A3(n99), .A4(n98), .ZN(n107) );
  aoi22d1 U11076 ( .A1(images_bus[189]), .A2(n435), .B1(images_bus[191]), .B2(
        n425), .ZN(n105) );
  aoi22d1 U11077 ( .A1(images_bus[185]), .A2(n454), .B1(n4958), .B2(n444), 
        .ZN(n104) );
  aoi22d1 U11078 ( .A1(images_bus[188]), .A2(n473), .B1(n6179), .B2(n463), 
        .ZN(n103) );
  aoi22d1 U11079 ( .A1(images_bus[184]), .A2(n491), .B1(images_bus[186]), .B2(
        n481), .ZN(n102) );
  nd04d0 U11080 ( .A1(n105), .A2(n104), .A3(n103), .A4(n102), .ZN(n106) );
  aoi22d1 U11081 ( .A1(n107), .A2(n385), .B1(n106), .B2(n383), .ZN(n119) );
  aoi22d1 U11082 ( .A1(images_bus[141]), .A2(n435), .B1(images_bus[143]), .B2(
        n425), .ZN(n111) );
  aoi22d1 U11083 ( .A1(images_bus[137]), .A2(n454), .B1(images_bus[139]), .B2(
        n444), .ZN(n110) );
  aoi22d1 U11084 ( .A1(images_bus[140]), .A2(n473), .B1(images_bus[142]), .B2(
        n463), .ZN(n109) );
  aoi22d1 U11085 ( .A1(images_bus[136]), .A2(n491), .B1(n6871), .B2(n481), 
        .ZN(n108) );
  nd04d0 U11086 ( .A1(n111), .A2(n110), .A3(n109), .A4(n108), .ZN(n117) );
  aoi22d1 U11087 ( .A1(images_bus[157]), .A2(n435), .B1(images_bus[159]), .B2(
        n425), .ZN(n115) );
  aoi22d1 U11088 ( .A1(images_bus[153]), .A2(n454), .B1(images_bus[155]), .B2(
        n444), .ZN(n114) );
  aoi22d1 U11089 ( .A1(images_bus[156]), .A2(n473), .B1(images_bus[158]), .B2(
        n463), .ZN(n113) );
  aoi22d1 U11090 ( .A1(images_bus[152]), .A2(n491), .B1(images_bus[154]), .B2(
        n479), .ZN(n112) );
  nd04d0 U11091 ( .A1(n115), .A2(n114), .A3(n113), .A4(n112), .ZN(n116) );
  aoi22d1 U11092 ( .A1(n117), .A2(n404), .B1(n116), .B2(n402), .ZN(n118) );
  oaim21d1 U11093 ( .B1(n119), .B2(n118), .A(n955), .ZN(n120) );
  aon211d1 U11094 ( .C1(n122), .C2(n121), .B(n955), .A(n120), .ZN(n123) );
  aoi22d1 U11095 ( .A1(n124), .A2(N3180), .B1(n123), .B2(n507), .ZN(n217) );
  aoi22d1 U11096 ( .A1(images_bus[101]), .A2(n435), .B1(images_bus[103]), .B2(
        n425), .ZN(n128) );
  aoi22d1 U11097 ( .A1(images_bus[97]), .A2(n454), .B1(images_bus[99]), .B2(
        n444), .ZN(n127) );
  aoi22d1 U11098 ( .A1(images_bus[100]), .A2(n473), .B1(images_bus[102]), .B2(
        n463), .ZN(n126) );
  aoi22d1 U11099 ( .A1(images_bus[96]), .A2(n491), .B1(images_bus[98]), .B2(
        n478), .ZN(n125) );
  nd04d0 U11100 ( .A1(n128), .A2(n127), .A3(n126), .A4(n125), .ZN(n134) );
  aoi22d1 U11101 ( .A1(images_bus[117]), .A2(n435), .B1(images_bus[119]), .B2(
        n425), .ZN(n132) );
  aoi22d1 U11102 ( .A1(images_bus[113]), .A2(n454), .B1(images_bus[115]), .B2(
        n444), .ZN(n131) );
  aoi22d1 U11103 ( .A1(n6547), .A2(n473), .B1(images_bus[118]), .B2(n463), 
        .ZN(n130) );
  aoi22d1 U11104 ( .A1(images_bus[112]), .A2(n491), .B1(n6795), .B2(n480), 
        .ZN(n129) );
  nd04d0 U11105 ( .A1(n132), .A2(n131), .A3(n130), .A4(n129), .ZN(n133) );
  aoi22d1 U11106 ( .A1(n134), .A2(n385), .B1(n133), .B2(n383), .ZN(n169) );
  aoi22d1 U11107 ( .A1(images_bus[69]), .A2(n434), .B1(images_bus[71]), .B2(
        n424), .ZN(n138) );
  aoi22d1 U11108 ( .A1(images_bus[65]), .A2(n453), .B1(images_bus[67]), .B2(
        n443), .ZN(n137) );
  aoi22d1 U11109 ( .A1(images_bus[68]), .A2(n472), .B1(images_bus[70]), .B2(
        n462), .ZN(n136) );
  aoi22d1 U11110 ( .A1(images_bus[64]), .A2(n490), .B1(images_bus[66]), .B2(
        n480), .ZN(n135) );
  nd04d0 U11111 ( .A1(n138), .A2(n137), .A3(n136), .A4(n135), .ZN(n144) );
  aoi22d1 U11112 ( .A1(images_bus[85]), .A2(n434), .B1(images_bus[87]), .B2(
        n424), .ZN(n142) );
  aoi22d1 U11113 ( .A1(images_bus[81]), .A2(n453), .B1(images_bus[83]), .B2(
        n443), .ZN(n141) );
  aoi22d1 U11114 ( .A1(images_bus[84]), .A2(n472), .B1(images_bus[86]), .B2(
        n462), .ZN(n140) );
  aoi22d1 U11115 ( .A1(images_bus[80]), .A2(n490), .B1(images_bus[82]), .B2(
        n477), .ZN(n139) );
  nd04d0 U11116 ( .A1(n142), .A2(n141), .A3(n140), .A4(n139), .ZN(n143) );
  aoi22d1 U11117 ( .A1(n144), .A2(n404), .B1(n143), .B2(n402), .ZN(n168) );
  aoi22d1 U11118 ( .A1(images_bus[109]), .A2(n434), .B1(images_bus[111]), .B2(
        n424), .ZN(n148) );
  aoi22d1 U11119 ( .A1(images_bus[105]), .A2(n453), .B1(images_bus[107]), .B2(
        n443), .ZN(n147) );
  aoi22d1 U11120 ( .A1(images_bus[108]), .A2(n472), .B1(images_bus[110]), .B2(
        n462), .ZN(n146) );
  aoi22d1 U11121 ( .A1(images_bus[104]), .A2(n490), .B1(images_bus[106]), .B2(
        n481), .ZN(n145) );
  nd04d0 U11122 ( .A1(n148), .A2(n147), .A3(n146), .A4(n145), .ZN(n154) );
  aoi22d1 U11123 ( .A1(images_bus[125]), .A2(n434), .B1(images_bus[127]), .B2(
        n424), .ZN(n152) );
  aoi22d1 U11124 ( .A1(images_bus[121]), .A2(n453), .B1(images_bus[123]), .B2(
        n443), .ZN(n151) );
  aoi22d1 U11125 ( .A1(images_bus[124]), .A2(n472), .B1(images_bus[126]), .B2(
        n462), .ZN(n150) );
  aoi22d1 U11126 ( .A1(images_bus[120]), .A2(n490), .B1(images_bus[122]), .B2(
        n480), .ZN(n149) );
  nd04d0 U11127 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .ZN(n153) );
  aoi22d1 U11128 ( .A1(n154), .A2(n385), .B1(n153), .B2(n383), .ZN(n166) );
  aoi22d1 U11129 ( .A1(images_bus[77]), .A2(n434), .B1(images_bus[79]), .B2(
        n424), .ZN(n158) );
  aoi22d1 U11130 ( .A1(images_bus[73]), .A2(n453), .B1(images_bus[75]), .B2(
        n443), .ZN(n157) );
  aoi22d1 U11131 ( .A1(images_bus[76]), .A2(n472), .B1(images_bus[78]), .B2(
        n462), .ZN(n156) );
  aoi22d1 U11132 ( .A1(images_bus[72]), .A2(n490), .B1(images_bus[74]), .B2(
        n479), .ZN(n155) );
  nd04d0 U11133 ( .A1(n158), .A2(n157), .A3(n156), .A4(n155), .ZN(n164) );
  aoi22d1 U11134 ( .A1(images_bus[93]), .A2(n434), .B1(images_bus[95]), .B2(
        n424), .ZN(n162) );
  aoi22d1 U11135 ( .A1(images_bus[89]), .A2(n453), .B1(images_bus[91]), .B2(
        n443), .ZN(n161) );
  aoi22d1 U11136 ( .A1(n6496), .A2(n472), .B1(images_bus[94]), .B2(n462), .ZN(
        n160) );
  aoi22d1 U11137 ( .A1(images_bus[88]), .A2(n490), .B1(n6699), .B2(n479), .ZN(
        n159) );
  nd04d0 U11138 ( .A1(n162), .A2(n161), .A3(n160), .A4(n159), .ZN(n163) );
  aoi22d1 U11139 ( .A1(n164), .A2(n404), .B1(n163), .B2(n402), .ZN(n165) );
  oaim21d1 U11140 ( .B1(n166), .B2(n165), .A(n955), .ZN(n167) );
  aon211d1 U11141 ( .C1(n169), .C2(n168), .B(n955), .A(n167), .ZN(n215) );
  aoi22d1 U11142 ( .A1(images_bus[37]), .A2(n434), .B1(images_bus[39]), .B2(
        n424), .ZN(n173) );
  aoi22d1 U11143 ( .A1(images_bus[33]), .A2(n453), .B1(images_bus[35]), .B2(
        n443), .ZN(n172) );
  aoi22d1 U11144 ( .A1(images_bus[36]), .A2(n472), .B1(images_bus[38]), .B2(
        n462), .ZN(n171) );
  aoi22d1 U11145 ( .A1(images_bus[32]), .A2(n490), .B1(n6967), .B2(n479), .ZN(
        n170) );
  nd04d0 U11146 ( .A1(n173), .A2(n172), .A3(n171), .A4(n170), .ZN(n179) );
  aoi22d1 U11147 ( .A1(n4331), .A2(n434), .B1(images_bus[55]), .B2(n424), .ZN(
        n177) );
  aoi22d1 U11148 ( .A1(images_bus[49]), .A2(n453), .B1(images_bus[51]), .B2(
        n443), .ZN(n176) );
  aoi22d1 U11149 ( .A1(images_bus[52]), .A2(n472), .B1(images_bus[54]), .B2(
        n462), .ZN(n175) );
  aoi22d1 U11150 ( .A1(images_bus[48]), .A2(n490), .B1(n6806), .B2(n479), .ZN(
        n174) );
  nd04d0 U11151 ( .A1(n177), .A2(n176), .A3(n175), .A4(n174), .ZN(n178) );
  aoi22d1 U11152 ( .A1(n179), .A2(n385), .B1(n178), .B2(n383), .ZN(n213) );
  aoi22d1 U11153 ( .A1(images_bus[5]), .A2(n434), .B1(images_bus[7]), .B2(n424), .ZN(n182) );
  aoi22d1 U11154 ( .A1(images_bus[1]), .A2(n453), .B1(images_bus[3]), .B2(n443), .ZN(n181) );
  aoi22d1 U11155 ( .A1(images_bus[4]), .A2(n472), .B1(images_bus[6]), .B2(n462), .ZN(n180) );
  nd04d0 U11156 ( .A1(n182), .A2(n181), .A3(n180), .A4(n3), .ZN(n188) );
  aoi22d1 U11157 ( .A1(images_bus[21]), .A2(n433), .B1(images_bus[23]), .B2(
        n423), .ZN(n186) );
  aoi22d1 U11158 ( .A1(images_bus[17]), .A2(n452), .B1(images_bus[19]), .B2(
        n442), .ZN(n185) );
  aoi22d1 U11159 ( .A1(images_bus[20]), .A2(n471), .B1(images_bus[22]), .B2(
        n461), .ZN(n184) );
  aoi22d1 U11160 ( .A1(images_bus[16]), .A2(n490), .B1(images_bus[18]), .B2(
        n479), .ZN(n183) );
  nd04d0 U11161 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(n187) );
  aoi22d1 U11162 ( .A1(n188), .A2(n404), .B1(n187), .B2(n402), .ZN(n212) );
  aoi22d1 U11163 ( .A1(images_bus[45]), .A2(n433), .B1(images_bus[47]), .B2(
        n423), .ZN(n192) );
  aoi22d1 U11164 ( .A1(images_bus[41]), .A2(n452), .B1(images_bus[43]), .B2(
        n442), .ZN(n191) );
  aoi22d1 U11165 ( .A1(images_bus[44]), .A2(n471), .B1(images_bus[46]), .B2(
        n461), .ZN(n190) );
  aoi22d1 U11166 ( .A1(images_bus[40]), .A2(n489), .B1(images_bus[42]), .B2(
        n479), .ZN(n189) );
  nd04d0 U11167 ( .A1(n192), .A2(n191), .A3(n190), .A4(n189), .ZN(n198) );
  aoi22d1 U11168 ( .A1(images_bus[61]), .A2(n433), .B1(images_bus[63]), .B2(
        n423), .ZN(n196) );
  aoi22d1 U11169 ( .A1(images_bus[57]), .A2(n452), .B1(images_bus[59]), .B2(
        n442), .ZN(n195) );
  aoi22d1 U11170 ( .A1(images_bus[60]), .A2(n471), .B1(images_bus[62]), .B2(
        n461), .ZN(n194) );
  aoi22d1 U11171 ( .A1(images_bus[56]), .A2(n489), .B1(images_bus[58]), .B2(
        n479), .ZN(n193) );
  nd04d0 U11172 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .ZN(n197) );
  aoi22d1 U11173 ( .A1(n198), .A2(n385), .B1(n197), .B2(n383), .ZN(n210) );
  aoi22d1 U11174 ( .A1(images_bus[13]), .A2(n433), .B1(images_bus[15]), .B2(
        n423), .ZN(n202) );
  aoi22d1 U11175 ( .A1(n5714), .A2(n452), .B1(images_bus[11]), .B2(n442), .ZN(
        n201) );
  aoi22d1 U11176 ( .A1(images_bus[12]), .A2(n471), .B1(images_bus[14]), .B2(
        n461), .ZN(n200) );
  aoi22d1 U11177 ( .A1(images_bus[8]), .A2(n489), .B1(n6890), .B2(n479), .ZN(
        n199) );
  nd04d0 U11178 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(n208) );
  aoi22d1 U11179 ( .A1(images_bus[29]), .A2(n433), .B1(images_bus[31]), .B2(
        n423), .ZN(n206) );
  aoi22d1 U11180 ( .A1(images_bus[25]), .A2(n452), .B1(images_bus[27]), .B2(
        n442), .ZN(n205) );
  aoi22d1 U11181 ( .A1(images_bus[28]), .A2(n471), .B1(images_bus[30]), .B2(
        n461), .ZN(n204) );
  aoi22d1 U11182 ( .A1(images_bus[24]), .A2(n489), .B1(images_bus[26]), .B2(
        n479), .ZN(n203) );
  nd04d0 U11183 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(n207) );
  aoi22d1 U11184 ( .A1(n208), .A2(n404), .B1(n207), .B2(n402), .ZN(n209) );
  oaim21d1 U11185 ( .B1(n210), .B2(n209), .A(n955), .ZN(n211) );
  aon211d1 U11186 ( .C1(n213), .C2(n212), .B(n955), .A(n211), .ZN(n214) );
  aoi22d1 U11187 ( .A1(n215), .A2(N3180), .B1(n214), .B2(n507), .ZN(n216) );
  oai22d1 U11188 ( .A1(n418), .A2(n217), .B1(N3181), .B2(n216), .ZN(n416) );
  aoi22d1 U11189 ( .A1(images_bus[485]), .A2(n433), .B1(images_bus[487]), .B2(
        n423), .ZN(n221) );
  aoi22d1 U11190 ( .A1(images_bus[481]), .A2(n452), .B1(images_bus[483]), .B2(
        n442), .ZN(n220) );
  aoi22d1 U11191 ( .A1(images_bus[484]), .A2(n471), .B1(images_bus[486]), .B2(
        n461), .ZN(n219) );
  aoi22d1 U11192 ( .A1(images_bus[480]), .A2(n489), .B1(n6892), .B2(n479), 
        .ZN(n218) );
  nd04d0 U11193 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(n227) );
  aoi22d1 U11194 ( .A1(n4297), .A2(n433), .B1(images_bus[503]), .B2(n423), 
        .ZN(n225) );
  aoi22d1 U11195 ( .A1(images_bus[497]), .A2(n452), .B1(images_bus[499]), .B2(
        n442), .ZN(n224) );
  aoi22d1 U11196 ( .A1(images_bus[500]), .A2(n471), .B1(images_bus[502]), .B2(
        n461), .ZN(n223) );
  aoi22d1 U11197 ( .A1(images_bus[496]), .A2(n489), .B1(images_bus[498]), .B2(
        n479), .ZN(n222) );
  nd04d0 U11198 ( .A1(n225), .A2(n224), .A3(n223), .A4(n222), .ZN(n226) );
  aoi22d1 U11199 ( .A1(n227), .A2(n385), .B1(n226), .B2(n383), .ZN(n262) );
  aoi22d1 U11200 ( .A1(images_bus[453]), .A2(n433), .B1(images_bus[455]), .B2(
        n423), .ZN(n231) );
  aoi22d1 U11201 ( .A1(images_bus[449]), .A2(n452), .B1(images_bus[451]), .B2(
        n442), .ZN(n230) );
  aoi22d1 U11202 ( .A1(n6598), .A2(n471), .B1(images_bus[454]), .B2(n461), 
        .ZN(n229) );
  aoi22d1 U11203 ( .A1(images_bus[448]), .A2(n489), .B1(images_bus[450]), .B2(
        n479), .ZN(n228) );
  nd04d0 U11204 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(n237) );
  aoi22d1 U11205 ( .A1(images_bus[469]), .A2(n433), .B1(images_bus[471]), .B2(
        n423), .ZN(n235) );
  aoi22d1 U11206 ( .A1(images_bus[465]), .A2(n452), .B1(images_bus[467]), .B2(
        n442), .ZN(n234) );
  aoi22d1 U11207 ( .A1(n6512), .A2(n471), .B1(n6212), .B2(n461), .ZN(n233) );
  aoi22d1 U11208 ( .A1(images_bus[464]), .A2(n489), .B1(images_bus[466]), .B2(
        n479), .ZN(n232) );
  nd04d0 U11209 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(n236) );
  aoi22d1 U11210 ( .A1(n237), .A2(n404), .B1(n236), .B2(n402), .ZN(n261) );
  aoi22d1 U11211 ( .A1(images_bus[493]), .A2(n432), .B1(images_bus[495]), .B2(
        n422), .ZN(n241) );
  aoi22d1 U11212 ( .A1(n5604), .A2(n451), .B1(images_bus[491]), .B2(n441), 
        .ZN(n240) );
  aoi22d1 U11213 ( .A1(images_bus[492]), .A2(n470), .B1(images_bus[494]), .B2(
        n460), .ZN(n239) );
  aoi22d1 U11214 ( .A1(images_bus[488]), .A2(n489), .B1(images_bus[490]), .B2(
        n478), .ZN(n238) );
  nd04d0 U11215 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(n247) );
  aoi22d1 U11216 ( .A1(images_bus[509]), .A2(n432), .B1(n6147), .B2(n422), 
        .ZN(n245) );
  aoi22d1 U11217 ( .A1(images_bus[505]), .A2(n451), .B1(images_bus[507]), .B2(
        n441), .ZN(n244) );
  aoi22d1 U11218 ( .A1(n6423), .A2(n470), .B1(n6152), .B2(n460), .ZN(n243) );
  aoi22d1 U11219 ( .A1(images_bus[504]), .A2(n488), .B1(images_bus[506]), .B2(
        n478), .ZN(n242) );
  nd04d0 U11220 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .ZN(n246) );
  aoi22d1 U11221 ( .A1(n247), .A2(n385), .B1(n246), .B2(n383), .ZN(n259) );
  aoi22d1 U11222 ( .A1(images_bus[461]), .A2(n432), .B1(images_bus[463]), .B2(
        n422), .ZN(n251) );
  aoi22d1 U11223 ( .A1(images_bus[457]), .A2(n451), .B1(images_bus[459]), .B2(
        n441), .ZN(n250) );
  aoi22d1 U11224 ( .A1(images_bus[460]), .A2(n470), .B1(n6279), .B2(n460), 
        .ZN(n249) );
  aoi22d1 U11225 ( .A1(images_bus[456]), .A2(n488), .B1(n6818), .B2(n478), 
        .ZN(n248) );
  nd04d0 U11226 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(n257) );
  aoi22d1 U11227 ( .A1(images_bus[477]), .A2(n432), .B1(images_bus[479]), .B2(
        n422), .ZN(n255) );
  aoi22d1 U11228 ( .A1(images_bus[473]), .A2(n451), .B1(images_bus[475]), .B2(
        n441), .ZN(n254) );
  aoi22d1 U11229 ( .A1(n6425), .A2(n470), .B1(n6155), .B2(n460), .ZN(n253) );
  aoi22d1 U11230 ( .A1(images_bus[472]), .A2(n488), .B1(images_bus[474]), .B2(
        n478), .ZN(n252) );
  nd04d0 U11231 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(n256) );
  aoi22d1 U11232 ( .A1(n257), .A2(n404), .B1(n256), .B2(n402), .ZN(n258) );
  oaim21d1 U11233 ( .B1(n259), .B2(n258), .A(n955), .ZN(n260) );
  aon211d1 U11234 ( .C1(n262), .C2(n261), .B(n955), .A(n260), .ZN(n309) );
  aoi22d1 U11235 ( .A1(images_bus[421]), .A2(n432), .B1(images_bus[423]), .B2(
        n422), .ZN(n266) );
  aoi22d1 U11236 ( .A1(images_bus[417]), .A2(n451), .B1(images_bus[419]), .B2(
        n441), .ZN(n265) );
  aoi22d1 U11237 ( .A1(n6599), .A2(n470), .B1(images_bus[422]), .B2(n460), 
        .ZN(n264) );
  aoi22d1 U11238 ( .A1(images_bus[416]), .A2(n488), .B1(images_bus[418]), .B2(
        n478), .ZN(n263) );
  nd04d0 U11239 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(n272) );
  aoi22d1 U11240 ( .A1(images_bus[437]), .A2(n432), .B1(images_bus[439]), .B2(
        n422), .ZN(n270) );
  aoi22d1 U11241 ( .A1(images_bus[433]), .A2(n451), .B1(images_bus[435]), .B2(
        n441), .ZN(n269) );
  aoi22d1 U11242 ( .A1(images_bus[436]), .A2(n470), .B1(images_bus[438]), .B2(
        n460), .ZN(n268) );
  aoi22d1 U11243 ( .A1(n7062), .A2(n488), .B1(images_bus[434]), .B2(n478), 
        .ZN(n267) );
  nd04d0 U11244 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(n271) );
  aoi22d1 U11245 ( .A1(n272), .A2(n385), .B1(n271), .B2(n383), .ZN(n307) );
  aoi22d1 U11246 ( .A1(images_bus[389]), .A2(n432), .B1(images_bus[391]), .B2(
        n422), .ZN(n276) );
  aoi22d1 U11247 ( .A1(images_bus[385]), .A2(n451), .B1(images_bus[387]), .B2(
        n441), .ZN(n275) );
  aoi22d1 U11248 ( .A1(n6600), .A2(n470), .B1(images_bus[390]), .B2(n460), 
        .ZN(n274) );
  aoi22d1 U11249 ( .A1(images_bus[384]), .A2(n488), .B1(n6901), .B2(n478), 
        .ZN(n273) );
  nd04d0 U11250 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .ZN(n282) );
  aoi22d1 U11251 ( .A1(images_bus[405]), .A2(n432), .B1(images_bus[407]), .B2(
        n422), .ZN(n280) );
  aoi22d1 U11252 ( .A1(images_bus[401]), .A2(n451), .B1(images_bus[403]), .B2(
        n441), .ZN(n279) );
  aoi22d1 U11253 ( .A1(images_bus[404]), .A2(n470), .B1(images_bus[406]), .B2(
        n460), .ZN(n278) );
  aoi22d1 U11254 ( .A1(images_bus[400]), .A2(n488), .B1(images_bus[402]), .B2(
        n478), .ZN(n277) );
  nd04d0 U11255 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(n281) );
  aoi22d1 U11256 ( .A1(n282), .A2(n404), .B1(n281), .B2(n402), .ZN(n306) );
  aoi22d1 U11257 ( .A1(images_bus[429]), .A2(n432), .B1(images_bus[431]), .B2(
        n422), .ZN(n286) );
  aoi22d1 U11258 ( .A1(images_bus[425]), .A2(n451), .B1(images_bus[427]), .B2(
        n441), .ZN(n285) );
  aoi22d1 U11259 ( .A1(n6556), .A2(n470), .B1(images_bus[430]), .B2(n460), 
        .ZN(n284) );
  aoi22d1 U11260 ( .A1(images_bus[424]), .A2(n488), .B1(images_bus[426]), .B2(
        n478), .ZN(n283) );
  nd04d0 U11261 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(n292) );
  aoi22d1 U11262 ( .A1(images_bus[445]), .A2(n431), .B1(images_bus[447]), .B2(
        n421), .ZN(n290) );
  aoi22d1 U11263 ( .A1(n5354), .A2(n450), .B1(images_bus[443]), .B2(n440), 
        .ZN(n289) );
  aoi22d1 U11264 ( .A1(images_bus[444]), .A2(n469), .B1(n6157), .B2(n459), 
        .ZN(n288) );
  aoi22d1 U11265 ( .A1(images_bus[440]), .A2(n488), .B1(images_bus[442]), .B2(
        n478), .ZN(n287) );
  nd04d0 U11266 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(n291) );
  aoi22d1 U11267 ( .A1(n385), .A2(n292), .B1(n383), .B2(n291), .ZN(n304) );
  aoi22d1 U11268 ( .A1(n4416), .A2(n431), .B1(images_bus[399]), .B2(n421), 
        .ZN(n296) );
  aoi22d1 U11269 ( .A1(images_bus[393]), .A2(n450), .B1(images_bus[395]), .B2(
        n440), .ZN(n295) );
  aoi22d1 U11270 ( .A1(images_bus[396]), .A2(n469), .B1(images_bus[398]), .B2(
        n459), .ZN(n294) );
  aoi22d1 U11271 ( .A1(images_bus[392]), .A2(n487), .B1(images_bus[394]), .B2(
        n478), .ZN(n293) );
  nd04d0 U11272 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(n302) );
  aoi22d1 U11273 ( .A1(images_bus[413]), .A2(n431), .B1(images_bus[415]), .B2(
        n421), .ZN(n300) );
  aoi22d1 U11274 ( .A1(images_bus[409]), .A2(n450), .B1(images_bus[411]), .B2(
        n440), .ZN(n299) );
  aoi22d1 U11275 ( .A1(n6437), .A2(n469), .B1(images_bus[414]), .B2(n459), 
        .ZN(n298) );
  aoi22d1 U11276 ( .A1(images_bus[408]), .A2(n487), .B1(n6659), .B2(n478), 
        .ZN(n297) );
  nd04d0 U11277 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .ZN(n301) );
  aoi22d1 U11278 ( .A1(n404), .A2(n302), .B1(n402), .B2(n301), .ZN(n303) );
  oaim21d1 U11279 ( .B1(n304), .B2(n303), .A(n955), .ZN(n305) );
  aon211d1 U11280 ( .C1(n307), .C2(n306), .B(n955), .A(n305), .ZN(n308) );
  aoi22d1 U11281 ( .A1(N3180), .A2(n309), .B1(n308), .B2(n507), .ZN(n414) );
  aoi22d1 U11282 ( .A1(images_bus[357]), .A2(n431), .B1(images_bus[359]), .B2(
        n421), .ZN(n313) );
  aoi22d1 U11283 ( .A1(images_bus[353]), .A2(n450), .B1(images_bus[355]), .B2(
        n440), .ZN(n312) );
  aoi22d1 U11284 ( .A1(n6601), .A2(n469), .B1(images_bus[358]), .B2(n459), 
        .ZN(n311) );
  aoi22d1 U11285 ( .A1(images_bus[352]), .A2(n487), .B1(n6908), .B2(n397), 
        .ZN(n310) );
  nd04d0 U11286 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(n319) );
  aoi22d1 U11287 ( .A1(images_bus[373]), .A2(n431), .B1(images_bus[375]), .B2(
        n421), .ZN(n317) );
  aoi22d1 U11288 ( .A1(images_bus[369]), .A2(n450), .B1(images_bus[371]), .B2(
        n440), .ZN(n316) );
  aoi22d1 U11289 ( .A1(images_bus[372]), .A2(n469), .B1(images_bus[374]), .B2(
        n459), .ZN(n315) );
  aoi22d1 U11290 ( .A1(images_bus[368]), .A2(n487), .B1(n6737), .B2(n397), 
        .ZN(n314) );
  nd04d0 U11291 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n318) );
  aoi22d1 U11292 ( .A1(n319), .A2(n385), .B1(n318), .B2(n383), .ZN(n354) );
  aoi22d1 U11293 ( .A1(images_bus[325]), .A2(n431), .B1(images_bus[327]), .B2(
        n421), .ZN(n323) );
  aoi22d1 U11294 ( .A1(images_bus[321]), .A2(n450), .B1(images_bus[323]), .B2(
        n440), .ZN(n322) );
  aoi22d1 U11295 ( .A1(images_bus[324]), .A2(n469), .B1(images_bus[326]), .B2(
        n459), .ZN(n321) );
  aoi22d1 U11296 ( .A1(images_bus[320]), .A2(n487), .B1(images_bus[322]), .B2(
        n480), .ZN(n320) );
  nd04d0 U11297 ( .A1(n323), .A2(n322), .A3(n321), .A4(n320), .ZN(n329) );
  aoi22d1 U11298 ( .A1(images_bus[341]), .A2(n431), .B1(images_bus[343]), .B2(
        n421), .ZN(n327) );
  aoi22d1 U11299 ( .A1(images_bus[337]), .A2(n450), .B1(images_bus[339]), .B2(
        n440), .ZN(n326) );
  aoi22d1 U11300 ( .A1(images_bus[340]), .A2(n469), .B1(n6235), .B2(n459), 
        .ZN(n325) );
  aoi22d1 U11301 ( .A1(images_bus[336]), .A2(n487), .B1(images_bus[338]), .B2(
        n397), .ZN(n324) );
  nd04d0 U11302 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(n328) );
  aoi22d1 U11303 ( .A1(n329), .A2(n404), .B1(n328), .B2(n402), .ZN(n353) );
  aoi22d1 U11304 ( .A1(images_bus[365]), .A2(n431), .B1(images_bus[367]), .B2(
        n421), .ZN(n333) );
  aoi22d1 U11305 ( .A1(n5626), .A2(n450), .B1(images_bus[363]), .B2(n440), 
        .ZN(n332) );
  aoi22d1 U11306 ( .A1(images_bus[364]), .A2(n469), .B1(images_bus[366]), .B2(
        n459), .ZN(n331) );
  aoi22d1 U11307 ( .A1(images_bus[360]), .A2(n487), .B1(images_bus[362]), .B2(
        n480), .ZN(n330) );
  nd04d0 U11308 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(n339) );
  aoi22d1 U11309 ( .A1(images_bus[381]), .A2(n431), .B1(images_bus[383]), .B2(
        n421), .ZN(n337) );
  aoi22d1 U11310 ( .A1(images_bus[377]), .A2(n450), .B1(images_bus[379]), .B2(
        n440), .ZN(n336) );
  aoi22d1 U11311 ( .A1(images_bus[380]), .A2(n469), .B1(images_bus[382]), .B2(
        n459), .ZN(n335) );
  aoi22d1 U11312 ( .A1(images_bus[376]), .A2(n487), .B1(n6664), .B2(n477), 
        .ZN(n334) );
  nd04d0 U11313 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .ZN(n338) );
  aoi22d1 U11314 ( .A1(n339), .A2(n385), .B1(n338), .B2(n383), .ZN(n351) );
  aoi22d1 U11315 ( .A1(images_bus[333]), .A2(n430), .B1(images_bus[335]), .B2(
        n420), .ZN(n343) );
  aoi22d1 U11316 ( .A1(images_bus[329]), .A2(n449), .B1(images_bus[331]), .B2(
        n439), .ZN(n342) );
  aoi22d1 U11317 ( .A1(images_bus[332]), .A2(n468), .B1(images_bus[334]), .B2(
        n458), .ZN(n341) );
  aoi22d1 U11318 ( .A1(images_bus[328]), .A2(n487), .B1(images_bus[330]), .B2(
        n478), .ZN(n340) );
  nd04d0 U11319 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(n349) );
  aoi22d1 U11320 ( .A1(images_bus[349]), .A2(n430), .B1(images_bus[351]), .B2(
        n420), .ZN(n347) );
  aoi22d1 U11321 ( .A1(images_bus[345]), .A2(n449), .B1(images_bus[347]), .B2(
        n439), .ZN(n346) );
  aoi22d1 U11322 ( .A1(images_bus[348]), .A2(n468), .B1(images_bus[350]), .B2(
        n458), .ZN(n345) );
  aoi22d1 U11323 ( .A1(images_bus[344]), .A2(n486), .B1(images_bus[346]), .B2(
        n477), .ZN(n344) );
  nd04d0 U11324 ( .A1(n347), .A2(n346), .A3(n345), .A4(n344), .ZN(n348) );
  aoi22d1 U11325 ( .A1(n349), .A2(n404), .B1(n348), .B2(n402), .ZN(n350) );
  oaim21d1 U11326 ( .B1(n351), .B2(n350), .A(n955), .ZN(n352) );
  aon211d1 U11327 ( .C1(n354), .C2(n353), .B(n955), .A(n352), .ZN(n412) );
  aoi22d1 U11328 ( .A1(images_bus[293]), .A2(n430), .B1(images_bus[295]), .B2(
        n420), .ZN(n358) );
  aoi22d1 U11329 ( .A1(images_bus[289]), .A2(n449), .B1(images_bus[291]), .B2(
        n439), .ZN(n357) );
  aoi22d1 U11330 ( .A1(images_bus[292]), .A2(n468), .B1(n6383), .B2(n458), 
        .ZN(n356) );
  aoi22d1 U11331 ( .A1(images_bus[288]), .A2(n486), .B1(n6922), .B2(n397), 
        .ZN(n355) );
  nd04d0 U11332 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(n364) );
  aoi22d1 U11333 ( .A1(images_bus[309]), .A2(n430), .B1(images_bus[311]), .B2(
        n420), .ZN(n362) );
  aoi22d1 U11334 ( .A1(images_bus[305]), .A2(n449), .B1(images_bus[307]), .B2(
        n439), .ZN(n361) );
  aoi22d1 U11335 ( .A1(n6531), .A2(n468), .B1(images_bus[310]), .B2(n458), 
        .ZN(n360) );
  aoi22d1 U11336 ( .A1(images_bus[304]), .A2(n486), .B1(images_bus[306]), .B2(
        n480), .ZN(n359) );
  nd04d0 U11337 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(n363) );
  aoi22d1 U11338 ( .A1(n364), .A2(n385), .B1(n363), .B2(n383), .ZN(n410) );
  aoi22d1 U11339 ( .A1(images_bus[261]), .A2(n430), .B1(images_bus[263]), .B2(
        n420), .ZN(n368) );
  aoi22d1 U11340 ( .A1(images_bus[257]), .A2(n449), .B1(images_bus[259]), .B2(
        n439), .ZN(n367) );
  aoi22d1 U11341 ( .A1(images_bus[260]), .A2(n468), .B1(images_bus[262]), .B2(
        n458), .ZN(n366) );
  aoi22d1 U11342 ( .A1(images_bus[256]), .A2(n486), .B1(images_bus[258]), .B2(
        n397), .ZN(n365) );
  nd04d0 U11343 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .ZN(n374) );
  aoi22d1 U11344 ( .A1(images_bus[277]), .A2(n430), .B1(images_bus[279]), .B2(
        n420), .ZN(n372) );
  aoi22d1 U11345 ( .A1(images_bus[273]), .A2(n449), .B1(images_bus[275]), .B2(
        n439), .ZN(n371) );
  aoi22d1 U11346 ( .A1(images_bus[276]), .A2(n468), .B1(images_bus[278]), .B2(
        n458), .ZN(n370) );
  aoi22d1 U11347 ( .A1(images_bus[272]), .A2(n486), .B1(images_bus[274]), .B2(
        n479), .ZN(n369) );
  nd04d0 U11348 ( .A1(n372), .A2(n371), .A3(n370), .A4(n369), .ZN(n373) );
  aoi22d1 U11349 ( .A1(n374), .A2(n404), .B1(n373), .B2(n402), .ZN(n409) );
  aoi22d1 U11350 ( .A1(images_bus[301]), .A2(n430), .B1(images_bus[303]), .B2(
        n420), .ZN(n378) );
  aoi22d1 U11351 ( .A1(images_bus[297]), .A2(n449), .B1(images_bus[299]), .B2(
        n439), .ZN(n377) );
  aoi22d1 U11352 ( .A1(images_bus[300]), .A2(n468), .B1(images_bus[302]), .B2(
        n458), .ZN(n376) );
  aoi22d1 U11353 ( .A1(images_bus[296]), .A2(n486), .B1(images_bus[298]), .B2(
        n477), .ZN(n375) );
  nd04d0 U11354 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(n386) );
  aoi22d1 U11355 ( .A1(images_bus[317]), .A2(n430), .B1(images_bus[319]), .B2(
        n420), .ZN(n382) );
  aoi22d1 U11356 ( .A1(images_bus[313]), .A2(n449), .B1(images_bus[315]), .B2(
        n439), .ZN(n381) );
  aoi22d1 U11357 ( .A1(images_bus[316]), .A2(n468), .B1(images_bus[318]), .B2(
        n458), .ZN(n380) );
  aoi22d1 U11358 ( .A1(images_bus[312]), .A2(n486), .B1(images_bus[314]), .B2(
        n477), .ZN(n379) );
  nd04d0 U11359 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(n384) );
  aoi22d1 U11360 ( .A1(n386), .A2(n385), .B1(n384), .B2(n383), .ZN(n407) );
  aoi22d1 U11361 ( .A1(images_bus[269]), .A2(n430), .B1(images_bus[271]), .B2(
        n420), .ZN(n390) );
  aoi22d1 U11362 ( .A1(images_bus[265]), .A2(n449), .B1(images_bus[267]), .B2(
        n439), .ZN(n389) );
  aoi22d1 U11363 ( .A1(images_bus[268]), .A2(n468), .B1(images_bus[270]), .B2(
        n458), .ZN(n388) );
  aoi22d1 U11364 ( .A1(images_bus[264]), .A2(n486), .B1(images_bus[266]), .B2(
        n477), .ZN(n387) );
  nd04d0 U11365 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(n405) );
  aoi22d1 U11366 ( .A1(images_bus[285]), .A2(n438), .B1(images_bus[287]), .B2(
        n429), .ZN(n401) );
  aoi22d1 U11367 ( .A1(images_bus[281]), .A2(n457), .B1(n4946), .B2(n448), 
        .ZN(n400) );
  aoi22d1 U11368 ( .A1(n6466), .A2(n476), .B1(images_bus[286]), .B2(n467), 
        .ZN(n399) );
  aoi22d1 U11369 ( .A1(images_bus[280]), .A2(n486), .B1(images_bus[282]), .B2(
        n477), .ZN(n398) );
  nd04d0 U11370 ( .A1(n401), .A2(n400), .A3(n399), .A4(n398), .ZN(n403) );
  aoi22d1 U11371 ( .A1(n405), .A2(n404), .B1(n403), .B2(n402), .ZN(n406) );
  oaim21d1 U11372 ( .B1(n407), .B2(n406), .A(n955), .ZN(n408) );
  aon211d1 U11373 ( .C1(n410), .C2(n409), .B(n955), .A(n408), .ZN(n411) );
  aoi22d1 U11374 ( .A1(n412), .A2(N3180), .B1(n411), .B2(n507), .ZN(n413) );
  oai22d1 U11375 ( .A1(n414), .A2(n418), .B1(n509), .B2(n413), .ZN(n415) );
  aor22d1 U11376 ( .A1(n416), .A2(n419), .B1(N3182), .B2(n415), .Z(N5285) );
  xr02d1 U11377 ( .A1(\add_0_root_add_1_root_add_98_3/carry[11] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[11] ), .Z(N3887) );
  an02d0 U11378 ( .A1(\add_0_root_add_1_root_add_98_3/A[10] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[10] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[11] ) );
  xr02d1 U11379 ( .A1(\add_0_root_add_1_root_add_98_3/carry[10] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[10] ), .Z(N3886) );
  an02d0 U11380 ( .A1(\add_0_root_add_1_root_add_98_3/A[9] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[9] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[10] ) );
  xr02d1 U11381 ( .A1(\add_0_root_add_1_root_add_98_3/carry[9] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[9] ), .Z(N3885) );
  or02d0 U11382 ( .A1(\add_0_root_add_1_root_add_98_3/carry[8] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[8] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[9] ) );
  xn02d1 U11383 ( .A1(\add_0_root_add_1_root_add_98_3/A[8] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[8] ), .ZN(N3884) );
  an02d0 U11384 ( .A1(\add_0_root_add_1_root_add_98_3/A[7] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[7] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[8] ) );
  xr02d1 U11385 ( .A1(\add_0_root_add_1_root_add_98_3/carry[7] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[7] ), .Z(N3883) );
  an02d0 U11386 ( .A1(\add_0_root_add_1_root_add_98_3/A[6] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[6] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[7] ) );
  xr02d1 U11387 ( .A1(\add_0_root_add_1_root_add_98_3/carry[6] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[6] ), .Z(N3882) );
  an02d0 U11388 ( .A1(\add_0_root_add_1_root_add_98_3/A[5] ), .A2(
        \add_0_root_add_1_root_add_98_3/carry[5] ), .Z(
        \add_0_root_add_1_root_add_98_3/carry[6] ) );
  xr02d1 U11389 ( .A1(\add_0_root_add_1_root_add_98_3/carry[5] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[5] ), .Z(N3881) );
  an02d0 U11390 ( .A1(\add_0_root_add_1_root_add_98_3/A[3] ), .A2(N3855), .Z(
        \add_0_root_add_1_root_add_98_3/carry[4] ) );
  xr02d1 U11391 ( .A1(N3855), .A2(\add_0_root_add_1_root_add_98_3/A[3] ), .Z(
        N3879) );
  xr02d1 U11392 ( .A1(\add_1_root_add_89_2/carry[11] ), .A2(
        temp_new_reference[8]), .Z(N3239) );
  an02d0 U11393 ( .A1(temp_new_reference[7]), .A2(
        \add_1_root_add_89_2/carry[10] ), .Z(\add_1_root_add_89_2/carry[11] )
         );
  xr02d1 U11394 ( .A1(\add_1_root_add_89_2/carry[10] ), .A2(
        temp_new_reference[7]), .Z(N3238) );
  an02d0 U11395 ( .A1(temp_new_reference[6]), .A2(temp_new_reference[5]), .Z(
        \add_1_root_add_89_2/carry[10] ) );
  xr02d1 U11396 ( .A1(temp_new_reference[5]), .A2(temp_new_reference[6]), .Z(
        N3237) );
  xr02d1 U11397 ( .A1(\add_1_root_add_158_3/carry[11] ), .A2(N4013), .Z(N5111)
         );
  an02d0 U11398 ( .A1(N4012), .A2(\add_1_root_add_158_3/carry[10] ), .Z(
        \add_1_root_add_158_3/carry[11] ) );
  xr02d1 U11399 ( .A1(\add_1_root_add_158_3/carry[10] ), .A2(N4012), .Z(N5110)
         );
  an02d0 U11400 ( .A1(N4011), .A2(N4010), .Z(\add_1_root_add_158_3/carry[10] )
         );
  xr02d1 U11401 ( .A1(N4010), .A2(N4011), .Z(N5109) );
  xr02d1 U11402 ( .A1(\add_1_root_add_115_2/carry[11] ), .A2(n510), .Z(N4004)
         );
  an02d0 U11403 ( .A1(N3181), .A2(\add_1_root_add_115_2/carry[10] ), .Z(
        \add_1_root_add_115_2/carry[11] ) );
  xr02d1 U11404 ( .A1(\add_1_root_add_115_2/carry[10] ), .A2(N3181), .Z(N4003)
         );
  an02d0 U11405 ( .A1(n508), .A2(n506), .Z(\add_1_root_add_115_2/carry[10] )
         );
  xr02d1 U11406 ( .A1(N3179), .A2(n508), .Z(N4002) );
  xr02d1 U11407 ( .A1(\add_0_root_add_1_root_add_130_3/carry[11] ), .A2(n510), 
        .Z(N4696) );
  an02d0 U11408 ( .A1(N3181), .A2(\add_0_root_add_1_root_add_130_3/carry[10] ), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[11] ) );
  xr02d1 U11409 ( .A1(\add_0_root_add_1_root_add_130_3/carry[10] ), .A2(N3181), 
        .Z(N4695) );
  an02d0 U11410 ( .A1(n508), .A2(\add_0_root_add_1_root_add_130_3/carry[9] ), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[10] ) );
  xr02d1 U11411 ( .A1(\add_0_root_add_1_root_add_130_3/carry[9] ), .A2(N3180), 
        .Z(N4694) );
  or02d0 U11412 ( .A1(\add_0_root_add_1_root_add_130_3/carry[8] ), .A2(n506), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[9] ) );
  xn02d1 U11413 ( .A1(N3179), .A2(\add_0_root_add_1_root_add_130_3/carry[8] ), 
        .ZN(N4693) );
  an02d0 U11414 ( .A1(n504), .A2(\add_0_root_add_1_root_add_130_3/carry[7] ), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[8] ) );
  xr02d1 U11415 ( .A1(\add_0_root_add_1_root_add_130_3/carry[7] ), .A2(N3976), 
        .Z(N4692) );
  an02d0 U11416 ( .A1(n955), .A2(\add_0_root_add_1_root_add_130_3/carry[6] ), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[7] ) );
  xr02d1 U11417 ( .A1(\add_0_root_add_1_root_add_130_3/carry[6] ), .A2(n955), 
        .Z(N4691) );
  an02d0 U11418 ( .A1(n502), .A2(\add_0_root_add_1_root_add_130_3/carry[5] ), 
        .Z(\add_0_root_add_1_root_add_130_3/carry[6] ) );
  xr02d1 U11419 ( .A1(\add_0_root_add_1_root_add_130_3/carry[5] ), .A2(n502), 
        .Z(N4690) );
  an02d0 U11420 ( .A1(n513), .A2(N4664), .Z(
        \add_0_root_add_1_root_add_130_3/carry[4] ) );
  xr02d1 U11421 ( .A1(N4664), .A2(N3972), .Z(N4688) );
  xr02d1 U11422 ( .A1(\add_0_root_add_0_root_add_97_2/carry[11] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[11] ), .Z(N3851) );
  an02d0 U11423 ( .A1(\add_0_root_add_1_root_add_98_3/A[10] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[10] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[11] ) );
  xr02d1 U11424 ( .A1(\add_0_root_add_0_root_add_97_2/carry[10] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[10] ), .Z(N3850) );
  an02d0 U11425 ( .A1(\add_0_root_add_1_root_add_98_3/A[9] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[9] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[10] ) );
  xr02d1 U11426 ( .A1(\add_0_root_add_0_root_add_97_2/carry[9] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[9] ), .Z(N3849) );
  or02d0 U11427 ( .A1(\add_0_root_add_0_root_add_97_2/carry[8] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[8] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[9] ) );
  xn02d1 U11428 ( .A1(\add_0_root_add_1_root_add_98_3/A[8] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[8] ), .ZN(N3848) );
  an02d0 U11429 ( .A1(\add_0_root_add_1_root_add_98_3/A[7] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[7] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[8] ) );
  xr02d1 U11430 ( .A1(\add_0_root_add_0_root_add_97_2/carry[7] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[7] ), .Z(N3847) );
  an02d0 U11431 ( .A1(\add_0_root_add_1_root_add_98_3/A[6] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[6] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[7] ) );
  xr02d1 U11432 ( .A1(\add_0_root_add_0_root_add_97_2/carry[6] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[6] ), .Z(N3846) );
  an02d0 U11433 ( .A1(\add_0_root_add_1_root_add_98_3/A[5] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[5] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[6] ) );
  xr02d1 U11434 ( .A1(\add_0_root_add_0_root_add_97_2/carry[5] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[5] ), .Z(N3845) );
  an02d0 U11435 ( .A1(\add_0_root_add_1_root_add_98_3/A[4] ), .A2(
        \add_0_root_add_0_root_add_97_2/carry[4] ), .Z(
        \add_0_root_add_0_root_add_97_2/carry[5] ) );
  xr02d1 U11436 ( .A1(\add_0_root_add_0_root_add_97_2/carry[4] ), .A2(
        \add_0_root_add_1_root_add_98_3/A[4] ), .Z(N3844) );
  an02d0 U11437 ( .A1(\add_0_root_add_1_root_add_98_3/A[3] ), .A2(N3855), .Z(
        \add_0_root_add_0_root_add_97_2/carry[4] ) );
  xr02d1 U11438 ( .A1(N3855), .A2(\add_0_root_add_1_root_add_98_3/A[3] ), .Z(
        N3843) );
  xr02d1 U11439 ( .A1(\add_88_aco/carry[11] ), .A2(N29417), .Z(N3215) );
  an02d0 U11440 ( .A1(N29416), .A2(\add_88_aco/carry[10] ), .Z(
        \add_88_aco/carry[11] ) );
  xr02d1 U11441 ( .A1(\add_88_aco/carry[10] ), .A2(N29416), .Z(N3214) );
  an02d0 U11442 ( .A1(N29415), .A2(N29414), .Z(\add_88_aco/carry[10] ) );
  xr02d1 U11443 ( .A1(N29414), .A2(N29415), .Z(N3213) );
  xr02d1 U11444 ( .A1(\add_157_2/carry[11] ), .A2(N4013), .Z(N5078) );
  an02d0 U11445 ( .A1(N4012), .A2(\add_157_2/carry[10] ), .Z(
        \add_157_2/carry[11] ) );
  xr02d1 U11446 ( .A1(\add_157_2/carry[10] ), .A2(N4012), .Z(N5077) );
  an02d0 U11447 ( .A1(N4011), .A2(N4010), .Z(\add_157_2/carry[10] ) );
  xr02d1 U11448 ( .A1(N4010), .A2(N4011), .Z(N5076) );
  xr02d1 U11449 ( .A1(\add_114/carry[11] ), .A2(n510), .Z(N3980) );
  an02d0 U11450 ( .A1(N3181), .A2(\add_114/carry[10] ), .Z(\add_114/carry[11] ) );
  xr02d1 U11451 ( .A1(\add_114/carry[10] ), .A2(N3181), .Z(N3979) );
  an02d0 U11452 ( .A1(n508), .A2(n506), .Z(\add_114/carry[10] ) );
  xr02d1 U11453 ( .A1(N3179), .A2(n508), .Z(N3978) );
  xr02d1 U11454 ( .A1(n510), .A2(\add_0_root_add_0_root_add_129_2/carry[11] ), 
        .Z(N4660) );
  an02d0 U11455 ( .A1(\add_0_root_add_0_root_add_129_2/carry[10] ), .A2(N3181), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[11] ) );
  xr02d1 U11456 ( .A1(N3181), .A2(\add_0_root_add_0_root_add_129_2/carry[10] ), 
        .Z(N4659) );
  an02d0 U11457 ( .A1(\add_0_root_add_0_root_add_129_2/carry[9] ), .A2(n508), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[10] ) );
  xr02d1 U11458 ( .A1(N3180), .A2(\add_0_root_add_0_root_add_129_2/carry[9] ), 
        .Z(N4658) );
  or02d0 U11459 ( .A1(n506), .A2(\add_0_root_add_0_root_add_129_2/carry[8] ), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[9] ) );
  xn02d1 U11460 ( .A1(\add_0_root_add_0_root_add_129_2/carry[8] ), .A2(N3179), 
        .ZN(N4657) );
  an02d0 U11461 ( .A1(\add_0_root_add_0_root_add_129_2/carry[7] ), .A2(n504), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[8] ) );
  xr02d1 U11462 ( .A1(n504), .A2(\add_0_root_add_0_root_add_129_2/carry[7] ), 
        .Z(N4656) );
  an02d0 U11463 ( .A1(\add_0_root_add_0_root_add_129_2/carry[6] ), .A2(n955), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[7] ) );
  xr02d1 U11464 ( .A1(n955), .A2(\add_0_root_add_0_root_add_129_2/carry[6] ), 
        .Z(N4655) );
  an02d0 U11465 ( .A1(\add_0_root_add_0_root_add_129_2/carry[5] ), .A2(n502), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[6] ) );
  xr02d1 U11466 ( .A1(n502), .A2(\add_0_root_add_0_root_add_129_2/carry[5] ), 
        .Z(N4654) );
  an02d0 U11467 ( .A1(\add_0_root_add_0_root_add_129_2/carry[4] ), .A2(N3973), 
        .Z(\add_0_root_add_0_root_add_129_2/carry[5] ) );
  xr02d1 U11468 ( .A1(N3973), .A2(\add_0_root_add_0_root_add_129_2/carry[4] ), 
        .Z(N4653) );
  an02d0 U11469 ( .A1(N3855), .A2(n513), .Z(
        \add_0_root_add_0_root_add_129_2/carry[4] ) );
  xr02d1 U11470 ( .A1(n513), .A2(N3855), .Z(N4652) );
  xn02d1 U11471 ( .A1(n1335), .A2(\sub_183/carry[8] ), .ZN(N6875) );
  or02d0 U11472 ( .A1(\sub_183/carry[7] ), .A2(n1303), .Z(\sub_183/carry[8] )
         );
  xn02d1 U11473 ( .A1(n1277), .A2(\sub_183/carry[7] ), .ZN(N6874) );
  or02d0 U11474 ( .A1(\sub_183/carry[6] ), .A2(n1248), .Z(\sub_183/carry[7] )
         );
  xn02d1 U11475 ( .A1(n1230), .A2(\sub_183/carry[6] ), .ZN(N6873) );
  or02d0 U11476 ( .A1(\sub_183/carry[5] ), .A2(n1178), .Z(\sub_183/carry[6] )
         );
  xn02d1 U11477 ( .A1(n1190), .A2(\sub_183/carry[5] ), .ZN(N6872) );
  or02d0 U11478 ( .A1(\sub_183/carry[4] ), .A2(n1158), .Z(\sub_183/carry[5] )
         );
  xn02d1 U11479 ( .A1(n1153), .A2(\sub_183/carry[4] ), .ZN(N6871) );
  or02d0 U11480 ( .A1(\sub_183/carry[3] ), .A2(n1117), .Z(\sub_183/carry[4] )
         );
  xn02d1 U11481 ( .A1(n1099), .A2(\sub_183/carry[3] ), .ZN(N6870) );
  or02d0 U11482 ( .A1(n1027), .A2(n1080), .Z(\sub_183/carry[3] ) );
  xn02d1 U11483 ( .A1(n1042), .A2(n998), .ZN(N6869) );
  an02d0 U11484 ( .A1(N27499), .A2(N28066), .Z(
        \add_3_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11485 ( .A1(N28066), .A2(N27499), .Z(N28498) );
  an02d0 U11486 ( .A1(N28084), .A2(N27553), .Z(
        \add_5_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11487 ( .A1(N27553), .A2(N28084), .Z(N28066) );
  an02d0 U11488 ( .A1(N28138), .A2(N27625), .Z(
        \add_17_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11489 ( .A1(N27625), .A2(N28138), .Z(N27553) );
  an02d0 U11490 ( .A1(N27796), .A2(N27832), .Z(
        \add_32_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11491 ( .A1(N27832), .A2(N27796), .Z(N27625) );
  an02d0 U11492 ( .A1(N27301), .A2(N28282), .Z(
        \add_79_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11493 ( .A1(N28282), .A2(N27301), .Z(N27832) );
  an02d0 U11494 ( .A1(N28597), .A2(N28552), .Z(
        \add_72_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11495 ( .A1(N28552), .A2(N28597), .Z(N27796) );
  an02d0 U11496 ( .A1(N28228), .A2(N27841), .Z(
        \add_36_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11497 ( .A1(N27841), .A2(N28228), .Z(N28138) );
  an02d0 U11498 ( .A1(N28030), .A2(N28561), .Z(
        \add_80_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11499 ( .A1(N28561), .A2(N28030), .Z(N27841) );
  an02d0 U11500 ( .A1(N27346), .A2(N27472), .Z(
        \add_75_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11501 ( .A1(N27472), .A2(N27346), .Z(N28228) );
  an02d0 U11502 ( .A1(N28381), .A2(N27598), .Z(
        \add_12_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11503 ( .A1(N27598), .A2(N28381), .Z(N28084) );
  an02d0 U11504 ( .A1(N27724), .A2(N28165), .Z(
        \add_28_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11505 ( .A1(N28165), .A2(N27724), .Z(N27598) );
  an02d0 U11506 ( .A1(N27940), .A2(N27112), .Z(
        \add_46_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11507 ( .A1(N27112), .A2(N27940), .Z(N28165) );
  an02d0 U11508 ( .A1(N27229), .A2(N28048), .Z(
        \add_55_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11509 ( .A1(N28048), .A2(N27229), .Z(N27724) );
  an02d0 U11510 ( .A1(N28525), .A2(N28183), .Z(
        \add_26_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11511 ( .A1(N28183), .A2(N28525), .Z(N28381) );
  an02d0 U11512 ( .A1(N28345), .A2(N27130), .Z(
        \add_54_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11513 ( .A1(N27130), .A2(N28345), .Z(N28183) );
  an02d0 U11514 ( .A1(N28264), .A2(N28453), .Z(
        \add_49_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11515 ( .A1(N28453), .A2(N28264), .Z(N28525) );
  an02d0 U11516 ( .A1(N27535), .A2(N27544), .Z(
        \add_7_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11517 ( .A1(N27544), .A2(N27535), .Z(N27499) );
  an02d0 U11518 ( .A1(N28579), .A2(N28516), .Z(
        \add_16_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11519 ( .A1(N28516), .A2(N28579), .Z(N27544) );
  an02d0 U11520 ( .A1(N27778), .A2(N27787), .Z(
        \add_34_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11521 ( .A1(N27787), .A2(N27778), .Z(N28516) );
  an02d0 U11522 ( .A1(N28336), .A2(N27922), .Z(
        \add_70_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11523 ( .A1(N27922), .A2(N28336), .Z(N27787) );
  an02d0 U11524 ( .A1(N28462), .A2(N27202), .Z(
        \add_69_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11525 ( .A1(N27202), .A2(N28462), .Z(N27778) );
  an02d0 U11526 ( .A1(N27760), .A2(N28237), .Z(
        \add_33_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11527 ( .A1(N28237), .A2(N27760), .Z(N28579) );
  an02d0 U11528 ( .A1(N27175), .A2(N27400), .Z(
        \add_78_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11529 ( .A1(N27400), .A2(N27175), .Z(N28237) );
  an02d0 U11530 ( .A1(N27274), .A2(N28273), .Z(
        \add_62_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11531 ( .A1(N28273), .A2(N27274), .Z(N27760) );
  an02d0 U11532 ( .A1(N27607), .A2(N27571), .Z(
        \add_14_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11533 ( .A1(N27571), .A2(N27607), .Z(N27535) );
  an02d0 U11534 ( .A1(N27697), .A2(N28417), .Z(
        \add_22_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11535 ( .A1(N28417), .A2(N27697), .Z(N27571) );
  an02d0 U11536 ( .A1(N27877), .A2(N27238), .Z(
        \add_57_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11537 ( .A1(N27238), .A2(N27877), .Z(N28417) );
  an02d0 U11538 ( .A1(N27445), .A2(N27949), .Z(
        \add_48_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11539 ( .A1(N27949), .A2(N27445), .Z(N27697) );
  an02d0 U11540 ( .A1(N27742), .A2(N27679), .Z(
        \add_29_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11541 ( .A1(N27679), .A2(N27742), .Z(N27607) );
  an02d0 U11542 ( .A1(N27994), .A2(N27121), .Z(
        \add_45_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11543 ( .A1(N27121), .A2(N27994), .Z(N27679) );
  an02d0 U11544 ( .A1(N27328), .A2(N27382), .Z(
        \add_59_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11545 ( .A1(N27382), .A2(N27328), .Z(N27742) );
  an02d0 U11546 ( .A1(N28354), .A2(N28570), .Z(
        \add_1_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11547 ( .A1(N28570), .A2(N28354), .Z(N28606) );
  an02d0 U11548 ( .A1(N27490), .A2(N28075), .Z(
        \add_2_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11549 ( .A1(N28075), .A2(N27490), .Z(N28570) );
  an02d0 U11550 ( .A1(N28372), .A2(N28507), .Z(
        \add_8_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11551 ( .A1(N28507), .A2(N28372), .Z(N28075) );
  an02d0 U11552 ( .A1(N27643), .A2(N28120), .Z(
        \add_18_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11553 ( .A1(N28120), .A2(N27643), .Z(N28507) );
  an02d0 U11554 ( .A1(N28192), .A2(N27688), .Z(
        \add_27_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11555 ( .A1(N27688), .A2(N28192), .Z(N28120) );
  an02d0 U11556 ( .A1(N27976), .A2(N27913), .Z(
        \add_47_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11557 ( .A1(N27913), .A2(N27976), .Z(N27688) );
  an02d0 U11558 ( .A1(N27967), .A2(N27454), .Z(
        \add_58_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11559 ( .A1(N27454), .A2(N27967), .Z(N28192) );
  an02d0 U11560 ( .A1(N27805), .A2(N28588), .Z(
        \add_38_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11561 ( .A1(N28588), .A2(N27805), .Z(N27643) );
  an02d0 U11562 ( .A1(N27220), .A2(N27409), .Z(
        \add_65_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11563 ( .A1(N27409), .A2(N27220), .Z(N28588) );
  an02d0 U11564 ( .A1(N28057), .A2(N28012), .Z(
        \add_73_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11565 ( .A1(N28012), .A2(N28057), .Z(N27805) );
  an02d0 U11566 ( .A1(N27634), .A2(N27562), .Z(
        \add_19_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11567 ( .A1(N27562), .A2(N27634), .Z(N28372) );
  an02d0 U11568 ( .A1(N27751), .A2(N28426), .Z(
        \add_21_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11569 ( .A1(N28426), .A2(N27751), .Z(N27562) );
  an02d0 U11570 ( .A1(N27985), .A2(N28489), .Z(
        \add_67_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11571 ( .A1(N28489), .A2(N27985), .Z(N28426) );
  an02d0 U11572 ( .A1(N27427), .A2(N28327), .Z(
        \add_60_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11573 ( .A1(N28327), .A2(N27427), .Z(N27751) );
  an02d0 U11574 ( .A1(N27814), .A2(N28534), .Z(
        \add_37_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11575 ( .A1(N28534), .A2(N27814), .Z(N27634) );
  an02d0 U11576 ( .A1(N27184), .A2(N27364), .Z(
        \add_66_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11577 ( .A1(N27364), .A2(N27184), .Z(N28534) );
  an02d0 U11578 ( .A1(N27355), .A2(N27211), .Z(
        \add_76_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11579 ( .A1(N27211), .A2(N27355), .Z(N27814) );
  an02d0 U11580 ( .A1(N27526), .A2(N28093), .Z(
        \add_6_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11581 ( .A1(N28093), .A2(N27526), .Z(N27490) );
  an02d0 U11582 ( .A1(N27652), .A2(N28147), .Z(
        \add_15_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11583 ( .A1(N28147), .A2(N27652), .Z(N28093) );
  an02d0 U11584 ( .A1(N27823), .A2(N28615), .Z(
        \add_39_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11585 ( .A1(N28615), .A2(N27823), .Z(N28147) );
  an02d0 U11586 ( .A1(N27886), .A2(N27895), .Z(
        \add_64_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11587 ( .A1(N27895), .A2(N27886), .Z(N28615) );
  an02d0 U11588 ( .A1(N28003), .A2(N27337), .Z(
        \add_77_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11589 ( .A1(N27337), .A2(N28003), .Z(N27823) );
  an02d0 U11590 ( .A1(N28444), .A2(N28246), .Z(
        \add_40_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11591 ( .A1(N28246), .A2(N28444), .Z(N27652) );
  an02d0 U11592 ( .A1(N28021), .A2(N27256), .Z(
        \add_82_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11593 ( .A1(N27256), .A2(N28021), .Z(N28444) );
  an02d0 U11594 ( .A1(N28129), .A2(N28111), .Z(
        \add_13_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11595 ( .A1(N28111), .A2(N28129), .Z(N27526) );
  an02d0 U11596 ( .A1(N28408), .A2(N28435), .Z(
        \add_23_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11597 ( .A1(N28435), .A2(N28408), .Z(N28111) );
  an02d0 U11598 ( .A1(N27193), .A2(N28480), .Z(
        \add_74_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11599 ( .A1(N28480), .A2(N27193), .Z(N28435) );
  an02d0 U11600 ( .A1(N27265), .A2(N27958), .Z(
        \add_50_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11601 ( .A1(N27958), .A2(N27265), .Z(N28408) );
  an02d0 U11602 ( .A1(N28201), .A2(N28543), .Z(
        \add_30_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11603 ( .A1(N28543), .A2(N28201), .Z(N28129) );
  an02d0 U11604 ( .A1(N27904), .A2(N28291), .Z(
        \add_81_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11605 ( .A1(N28291), .A2(N27904), .Z(N28543) );
  an02d0 U11606 ( .A1(N28255), .A2(N27391), .Z(
        \add_61_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11607 ( .A1(N27391), .A2(N28255), .Z(N28201) );
  an02d0 U11608 ( .A1(\add_4_root_add_86_root_add_255_countones_143/carry[5] ), 
        .A2(N27513), .Z(N28360) );
  xr02d1 U11609 ( .A1(N27513), .A2(
        \add_4_root_add_86_root_add_255_countones_143/carry[5] ), .Z(N28359)
         );
  an02d0 U11610 ( .A1(N28363), .A2(N27508), .Z(
        \add_4_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11611 ( .A1(N27508), .A2(N28363), .Z(N28354) );
  an02d0 U11612 ( .A1(N27589), .A2(N27580), .Z(
        \add_11_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11613 ( .A1(N27580), .A2(N27589), .Z(N28363) );
  an02d0 U11614 ( .A1(N28174), .A2(N27733), .Z(
        \add_24_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11615 ( .A1(N27733), .A2(N28174), .Z(N27580) );
  an02d0 U11616 ( .A1(N27931), .A2(N28300), .Z(
        \add_56_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11617 ( .A1(N28300), .A2(N27931), .Z(N27733) );
  an02d0 U11618 ( .A1(N28471), .A2(N27463), .Z(
        \add_51_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11619 ( .A1(N27463), .A2(N28471), .Z(N28174) );
  an02d0 U11620 ( .A1(N27706), .A2(N27769), .Z(
        \add_25_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11621 ( .A1(N27769), .A2(N27706), .Z(N27589) );
  an02d0 U11622 ( .A1(N27418), .A2(N27373), .Z(
        \add_63_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11623 ( .A1(N27373), .A2(N27418), .Z(N27769) );
  an02d0 U11624 ( .A1(N28039), .A2(N27247), .Z(
        \add_52_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11625 ( .A1(N27247), .A2(N28039), .Z(N27706) );
  an02d0 U11626 ( .A1(N28102), .A2(N27517), .Z(
        \add_9_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11627 ( .A1(N27517), .A2(N28102), .Z(N27508) );
  an02d0 U11628 ( .A1(N27616), .A2(N28390), .Z(
        \add_10_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11629 ( .A1(N28390), .A2(N27616), .Z(N27517) );
  an02d0 U11630 ( .A1(N28219), .A2(N28210), .Z(
        \add_35_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11631 ( .A1(N28210), .A2(N28219), .Z(N28390) );
  an02d0 U11632 ( .A1(N27481), .A2(N27166), .Z(
        \add_68_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11633 ( .A1(N27166), .A2(N27481), .Z(N28210) );
  an02d0 U11634 ( .A1(N28309), .A2(N28318), .Z(
        \add_71_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11635 ( .A1(N28318), .A2(N28309), .Z(N28219) );
  an02d0 U11636 ( .A1(N28156), .A2(N27670), .Z(
        \add_31_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11637 ( .A1(N27670), .A2(N28156), .Z(N27616) );
  an02d0 U11638 ( .A1(N27868), .A2(N27148), .Z(
        \add_44_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11639 ( .A1(N27148), .A2(N27868), .Z(N27670) );
  an02d0 U11640 ( .A1(N27292), .A2(N27319), .Z(
        \add_43_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11641 ( .A1(N27319), .A2(N27292), .Z(N28156) );
  an02d0 U11642 ( .A1(\add_20_root_add_86_root_add_255_countones_143/carry[3] ), .A2(N27664), .Z(N28106) );
  xr02d1 U11643 ( .A1(N27664), .A2(
        \add_20_root_add_86_root_add_255_countones_143/carry[3] ), .Z(N28105)
         );
  an02d0 U11644 ( .A1(N27715), .A2(N27661), .Z(
        \add_20_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11645 ( .A1(N27661), .A2(N27715), .Z(N28102) );
  an02d0 U11646 ( .A1(N27310), .A2(N27139), .Z(
        \add_53_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11647 ( .A1(N27139), .A2(N27310), .Z(N27715) );
  an02d0 U11648 ( .A1(\add_41_root_add_86_root_add_255_countones_143/carry[2] ), .A2(N28401), .Z(N27664) );
  xr02d1 U11649 ( .A1(N28401), .A2(
        \add_41_root_add_86_root_add_255_countones_143/carry[2] ), .Z(N27663)
         );
  an02d0 U11650 ( .A1(N27436), .A2(N28399), .Z(
        \add_41_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11651 ( .A1(N28399), .A2(N27436), .Z(N27661) );
  an02d0 U11652 ( .A1(N27283), .A2(N27859), .Z(
        \add_42_root_add_86_root_add_255_countones_143/carry[1] ) );
  xr02d1 U11653 ( .A1(N27859), .A2(N27283), .Z(N28399) );
  an02d0 U11654 ( .A1(temp_new_reference[7]), .A2(N26489), .Z(N29416) );
  an02d0 U11655 ( .A1(temp_new_reference[8]), .A2(N26489), .Z(N29417) );
  an02d0 U11656 ( .A1(N3231), .A2(N26489), .Z(N3207) );
  an02d0 U11657 ( .A1(N3232), .A2(N26489), .Z(N3208) );
  an02d0 U11658 ( .A1(N3233), .A2(N26489), .Z(N3209) );
  an02d0 U11659 ( .A1(N3234), .A2(N26489), .Z(N3210) );
  an02d0 U11660 ( .A1(N3235), .A2(N26489), .Z(N3211) );
  an02d0 U11661 ( .A1(temp_new_reference[5]), .A2(N26489), .Z(N29414) );
  an02d0 U11662 ( .A1(N26489), .A2(temp_new_reference[6]), .Z(N29415) );
  an02d0 U11663 ( .A1(N3877), .A2(N26480), .Z(N29399) );
  an02d0 U11664 ( .A1(N3878), .A2(N26480), .Z(N29400) );
  an02d0 U11665 ( .A1(N26480), .A2(N3855), .Z(N29401) );
  an02d0 U11666 ( .A1(N3877), .A2(N26480), .Z(N29403) );
  an02d0 U11667 ( .A1(N3878), .A2(N26480), .Z(N29404) );
  an02d0 U11668 ( .A1(N26480), .A2(N3855), .Z(N29405) );
  nd12d0 U11669 ( .A1(n1027), .A2(n993), .ZN(n1373) );
  oaim21d1 U11670 ( .B1(n978), .B2(n1015), .A(n1373), .ZN(N5113) );
  or02d0 U11671 ( .A1(n1373), .A2(n1038), .Z(n1374) );
  oaim21d1 U11672 ( .B1(n1373), .B2(n1063), .A(n1374), .ZN(N5114) );
  or02d0 U11673 ( .A1(n1374), .A2(n1116), .Z(n1375) );
  oaim21d1 U11674 ( .B1(n1374), .B2(n1099), .A(n1375), .ZN(N5115) );
  or02d0 U11675 ( .A1(n1375), .A2(n1158), .Z(n1376) );
  oaim21d1 U11676 ( .B1(n1375), .B2(n1156), .A(n1376), .ZN(N5116) );
  or02d0 U11677 ( .A1(n1376), .A2(n1181), .Z(n1377) );
  oaim21d1 U11678 ( .B1(n1376), .B2(n1193), .A(n1377), .ZN(N5117) );
  nr02d0 U11679 ( .A1(n1377), .A2(n1250), .ZN(n1378) );
  oaim21d1 U11680 ( .B1(n1377), .B2(n1237), .A(n1380), .ZN(N5118) );
  xr02d1 U11681 ( .A1(n1292), .A2(n1378), .Z(N5119) );
  nr03d0 U11682 ( .A1(n1307), .A2(n1347), .A3(n1380), .ZN(N5121) );
  oan211d1 U11683 ( .C1(n1380), .C2(n1276), .B(n1326), .A(N5121), .ZN(n1379)
         );
  nd02d0 U11684 ( .A1(N5119), .A2(n418), .ZN(n1388) );
  oai21d1 U11685 ( .B1(n508), .B2(n1399), .A(n1388), .ZN(n1381) );
  aoi22d1 U11686 ( .A1(n499), .A2(N5113), .B1(n512), .B2(n993), .ZN(n1383) );
  nd02d0 U11687 ( .A1(N5115), .A2(n956), .ZN(n1386) );
  nd03d0 U11688 ( .A1(n1386), .A2(n1396), .A3(n502), .ZN(n1382) );
  oai21d1 U11689 ( .B1(N5115), .B2(n956), .A(n1382), .ZN(n1385) );
  aoim211d1 U11690 ( .C1(N5113), .C2(n499), .A(n1383), .B(n1385), .ZN(n1384)
         );
  oan211d1 U11691 ( .C1(n502), .C2(n1396), .B(n1386), .A(n1385), .ZN(n1387) );
  nr02d0 U11692 ( .A1(n1398), .A2(n506), .ZN(n1390) );
  aoim211d1 U11693 ( .C1(n1397), .C2(n504), .A(n1387), .B(n1390), .ZN(n1394)
         );
  nd03d0 U11694 ( .A1(n1388), .A2(n1399), .A3(n508), .ZN(n1389) );
  oai21d1 U11695 ( .B1(N5119), .B2(n418), .A(n1389), .ZN(n1392) );
  aoi321d1 U11696 ( .C1(n1401), .C2(n1397), .C3(n504), .B1(n506), .B2(n1398), 
        .A(n1392), .ZN(n1391) );
  aoim21d1 U11697 ( .B1(n1392), .B2(n1402), .A(n1391), .ZN(n1393) );
  aoi321d1 U11698 ( .C1(n1402), .C2(n1403), .C3(n1394), .B1(n510), .B2(n1400), 
        .A(n1393), .ZN(n1395) );
  aoim211d1 U11699 ( .C1(n1400), .C2(n510), .A(n1395), .B(N5121), .ZN(N5122)
         );
  or02d0 U11700 ( .A1(distance[5]), .A2(n12085), .Z(n1412) );
  an02d0 U11701 ( .A1(temp_minimum[3]), .A2(n12082), .Z(n1405) );
  nr03d0 U11702 ( .A1(n1405), .A2(temp_minimum[2]), .A3(n12080), .ZN(n1404) );
  aoim21d1 U11703 ( .B1(temp_minimum[3]), .B2(n12082), .A(n1404), .ZN(n1407)
         );
  aon211d1 U11704 ( .C1(temp_minimum[2]), .C2(n12080), .B(n1405), .A(n1407), 
        .ZN(n1406) );
  oai211d1 U11705 ( .C1(distance[4]), .C2(n12083), .A(n1412), .B(n1406), .ZN(
        n1417) );
  aoim22d1 U11706 ( .A1(temp_minimum[0]), .A2(n12076), .B1(n12077), .B2(
        distance[1]), .Z(n1408) );
  aoi211d1 U11707 ( .C1(distance[1]), .C2(n12077), .A(n1419), .B(n1408), .ZN(
        n1416) );
  nd02d0 U11708 ( .A1(temp_minimum[7]), .A2(n12090), .ZN(n1409) );
  oai21d1 U11709 ( .B1(distance[6]), .B2(n12087), .A(n1409), .ZN(n1415) );
  nd03d0 U11710 ( .A1(n1409), .A2(n12087), .A3(distance[6]), .ZN(n1410) );
  oai21d1 U11711 ( .B1(temp_minimum[7]), .B2(n12090), .A(n1410), .ZN(n1411) );
  aoi321d1 U11712 ( .C1(distance[4]), .C2(n12083), .C3(n1412), .B1(n12085), 
        .B2(distance[5]), .A(n1411), .ZN(n1413) );
  aor21d1 U11713 ( .B1(n1415), .B2(n1420), .A(n1413), .Z(n1414) );
  oai321d1 U11714 ( .C1(n1417), .C2(n1416), .C3(n1415), .B1(temp_minimum[8]), 
        .B2(n12092), .A(n1414), .ZN(n1418) );
  nd04d0 U11715 ( .A1(n1328), .A2(n1304), .A3(n1254), .A4(n1188), .ZN(n1423)
         );
  nd03d0 U11716 ( .A1(n1023), .A2(n983), .A3(n1073), .ZN(n1422) );
  nd02d0 U11717 ( .A1(n1161), .A2(n1090), .ZN(n1421) );
  nr03d0 U11718 ( .A1(n1423), .A2(n1422), .A3(n1421), .ZN(N15633) );
  nd04d0 U11719 ( .A1(n1162), .A2(n1094), .A3(n1083), .A4(n1023), .ZN(n1425)
         );
  nd04d0 U11720 ( .A1(n1327), .A2(n1294), .A3(n1254), .A4(n1187), .ZN(n1424)
         );
  nr02d0 U11721 ( .A1(n1425), .A2(n1424), .ZN(N15618) );
  nd04d0 U11722 ( .A1(N11556), .A2(n1274), .A3(n1254), .A4(n1191), .ZN(n1428)
         );
  oai21d1 U11723 ( .B1(n969), .B2(n1011), .A(n1061), .ZN(n1427) );
  nd02d0 U11724 ( .A1(n1161), .A2(n1116), .ZN(n1426) );
  nr03d0 U11725 ( .A1(n1428), .A2(n1427), .A3(n1426), .ZN(N15602) );
  nd04d0 U11726 ( .A1(n1195), .A2(n1143), .A3(n1104), .A4(n1071), .ZN(n1430)
         );
  nd03d0 U11727 ( .A1(num_images[7]), .A2(n1257), .A3(N11556), .ZN(n1429) );
  nr02d0 U11728 ( .A1(n1430), .A2(n1429), .ZN(N15586) );
  nd03d0 U11729 ( .A1(n1272), .A2(n1257), .A3(N11556), .ZN(n1433) );
  an03d0 U11730 ( .A1(n1022), .A2(n978), .A3(n1116), .Z(n1431) );
  aon211d1 U11731 ( .C1(n1047), .C2(n1089), .B(n1431), .A(n1142), .ZN(n1432)
         );
  nr13d1 U11732 ( .A1(n1204), .A2(n1433), .A3(n1432), .ZN(N15570) );
  nd03d0 U11733 ( .A1(n1297), .A2(n1256), .A3(N11556), .ZN(n1436) );
  oai21d1 U11734 ( .B1(n1013), .B2(n1058), .A(n1105), .ZN(n1435) );
  nd02d0 U11735 ( .A1(n1205), .A2(n1158), .ZN(n1434) );
  nr03d0 U11736 ( .A1(n1436), .A2(n1435), .A3(n1434), .ZN(N15554) );
  nd03d0 U11737 ( .A1(n1300), .A2(n1256), .A3(N11556), .ZN(n1439) );
  oai21d1 U11738 ( .B1(n970), .B2(n1011), .A(n1105), .ZN(n1437) );
  aon211d1 U11739 ( .C1(n1047), .C2(n1089), .B(n1440), .A(n1143), .ZN(n1438)
         );
  nr13d1 U11740 ( .A1(n1204), .A2(n1439), .A3(n1438), .ZN(N15538) );
  an03d0 U11741 ( .A1(n1161), .A2(n1116), .A3(n1186), .Z(n1441) );
  an04d0 U11742 ( .A1(n1305), .A2(n1244), .A3(n1340), .A4(n1441), .Z(N15522)
         );
  aor31d1 U11743 ( .B1(n1018), .B2(n976), .B3(n1052), .A(n1105), .Z(n1443) );
  an03d0 U11744 ( .A1(n1308), .A2(n1248), .A3(n1339), .Z(n1442) );
  nd03d0 U11745 ( .A1(n1298), .A2(n1256), .A3(N11556), .ZN(n1445) );
  aon211d1 U11746 ( .C1(n1047), .C2(num_images[1]), .B(n1090), .A(n1141), .ZN(
        n1444) );
  nr13d1 U11747 ( .A1(n1204), .A2(n1445), .A3(n1444), .ZN(N15490) );
  an02d0 U11748 ( .A1(n1201), .A2(n1155), .Z(n1446) );
  oai321d1 U11749 ( .C1(n965), .C2(n1100), .C3(n1007), .B1(n1090), .B2(n1063), 
        .A(n1446), .ZN(n1448) );
  nd03d0 U11750 ( .A1(n1292), .A2(n1256), .A3(N11556), .ZN(n1447) );
  nr02d0 U11751 ( .A1(n1448), .A2(n1447), .ZN(N15474) );
  oai211d1 U11752 ( .C1(n1042), .C2(n1120), .A(n1153), .B(n1189), .ZN(n1450)
         );
  nd03d0 U11753 ( .A1(n1273), .A2(n1257), .A3(n1338), .ZN(n1449) );
  nr02d0 U11754 ( .A1(n1450), .A2(n1449), .ZN(N15458) );
  nd03d0 U11755 ( .A1(n1279), .A2(n1256), .A3(n1339), .ZN(n1452) );
  aoi211d1 U11756 ( .C1(n1014), .C2(n967), .A(n1102), .B(n1045), .ZN(n1451) );
  nr04d0 U11757 ( .A1(n1452), .A2(n1210), .A3(n1451), .A4(n1171), .ZN(N15442)
         );
  ora311d1 U11758 ( .C1(n1108), .C2(n1044), .C3(n1028), .A(n1155), .B(n1196), 
        .Z(n1453) );
  nd03d0 U11759 ( .A1(n1295), .A2(n1256), .A3(n1336), .ZN(n1455) );
  nr04d0 U11760 ( .A1(n1117), .A2(n1070), .A3(n1027), .A4(n979), .ZN(n1454) );
  nr04d0 U11761 ( .A1(n1455), .A2(n1176), .A3(n1454), .A4(n1171), .ZN(N15410)
         );
  an03d0 U11762 ( .A1(n1204), .A2(n1157), .A3(n1246), .Z(n1456) );
  an03d0 U11763 ( .A1(n1344), .A2(n1301), .A3(n1456), .Z(N15394) );
  an04d0 U11764 ( .A1(n1091), .A2(n1077), .A3(n1020), .A4(n978), .Z(n1457) );
  ora211d1 U11765 ( .C1(n1141), .C2(n1457), .A(n1248), .B(n1295), .Z(n1458) );
  an03d0 U11766 ( .A1(n1344), .A2(n1180), .A3(n1458), .Z(N15378) );
  aor31d1 U11767 ( .B1(n1069), .B2(n1016), .B3(n1093), .A(n1147), .Z(n1459) );
  an03d0 U11768 ( .A1(n1204), .A2(n1459), .A3(n1246), .Z(n1460) );
  an03d0 U11769 ( .A1(n1344), .A2(n1301), .A3(n1460), .Z(N15362) );
  ora211d1 U11770 ( .C1(n963), .C2(n1013), .A(n1081), .B(n1112), .Z(n1461) );
  ora211d1 U11771 ( .C1(n1137), .C2(n1461), .A(n1228), .B(n1295), .Z(n1462) );
  an03d0 U11772 ( .A1(n1344), .A2(num_images[5]), .A3(n1462), .Z(N15346) );
  nd02d0 U11773 ( .A1(n1345), .A2(n1304), .ZN(n1464) );
  aon211d1 U11774 ( .C1(n1090), .C2(n1045), .B(n1153), .A(n1192), .ZN(n1463)
         );
  nr13d1 U11775 ( .A1(n1252), .A2(n1464), .A3(n1463), .ZN(N15330) );
  aoi321d1 U11776 ( .C1(n969), .C2(n1091), .C3(n1006), .B1(n1107), .B2(n1054), 
        .A(n1155), .ZN(n1465) );
  nr23d1 U11777 ( .A1(n1256), .A2(num_images[7]), .A3(n1465), .ZN(n1466) );
  an03d0 U11778 ( .A1(n1344), .A2(n1184), .A3(n1466), .Z(N15314) );
  oan211d1 U11779 ( .C1(n1007), .C2(n1047), .B(n1094), .A(n1140), .ZN(n1467)
         );
  nr23d1 U11780 ( .A1(n1208), .A2(n1227), .A3(n1467), .ZN(n1468) );
  an03d0 U11781 ( .A1(n1344), .A2(n1301), .A3(n1468), .Z(N15298) );
  aoi21d1 U11782 ( .B1(n1101), .B2(n1049), .A(n1149), .ZN(n1470) );
  oai21d1 U11783 ( .B1(n970), .B2(n1010), .A(n1104), .ZN(n1469) );
  aoi21d1 U11784 ( .B1(n1470), .B2(n1469), .A(n1268), .ZN(n1471) );
  an04d0 U11785 ( .A1(n1343), .A2(n1201), .A3(n1471), .A4(n1295), .Z(N15282)
         );
  ora211d1 U11786 ( .C1(n1090), .C2(n1145), .A(n1187), .B(n1241), .Z(n1472) );
  an03d0 U11787 ( .A1(n1344), .A2(n1301), .A3(n1472), .Z(N15266) );
  aor311d1 U11788 ( .C1(n1017), .C2(n976), .C3(n1050), .A(n1147), .B(n1100), 
        .Z(n1473) );
  an03d0 U11789 ( .A1(n1252), .A2(n1473), .A3(n1300), .Z(n1474) );
  an03d0 U11790 ( .A1(n1344), .A2(n1178), .A3(n1474), .Z(N15250) );
  aor211d1 U11791 ( .C1(n1067), .C2(n1006), .A(n1137), .B(n1094), .Z(n1475) );
  an03d0 U11792 ( .A1(n1204), .A2(n1248), .A3(n1475), .Z(n1476) );
  an03d0 U11793 ( .A1(n1344), .A2(n1301), .A3(n1476), .Z(N15234) );
  oai21d1 U11794 ( .B1(n971), .B2(n1011), .A(n1061), .ZN(n1477) );
  ora311d1 U11795 ( .C1(n1146), .C2(n1111), .C3(n1479), .A(n1244), .B(n1275), 
        .Z(n1478) );
  an03d0 U11796 ( .A1(n1344), .A2(n1186), .A3(n1478), .Z(N15218) );
  oai21d1 U11797 ( .B1(n1060), .B2(n1097), .A(n1201), .ZN(n1480) );
  oaim21d1 U11798 ( .B1(n1156), .B2(n1193), .A(n1480), .ZN(n1481) );
  an04d0 U11799 ( .A1(n1342), .A2(n1299), .A3(n1246), .A4(n1481), .Z(N15202)
         );
  aor21d1 U11800 ( .B1(n1018), .B2(n971), .A(n1061), .Z(n1482) );
  ora311d1 U11801 ( .C1(n1145), .C2(n1119), .C3(n1482), .A(n1229), .B(n1293), 
        .Z(n1483) );
  an03d0 U11802 ( .A1(n1344), .A2(n1177), .A3(n1483), .Z(N15186) );
  or04d0 U11803 ( .A1(n1136), .A2(n1112), .A3(n1067), .A4(n1014), .Z(n1484) );
  an03d0 U11804 ( .A1(n1204), .A2(n1247), .A3(n1484), .Z(n1485) );
  an03d0 U11805 ( .A1(n1344), .A2(n1274), .A3(n1485), .Z(N15170) );
  or03d0 U11806 ( .A1(num_images[4]), .A2(n1117), .A3(n1038), .Z(n1486) );
  ora311d1 U11807 ( .C1(n1001), .C2(n962), .C3(n1486), .A(n1244), .B(n1293), 
        .Z(n1487) );
  an03d0 U11808 ( .A1(n1344), .A2(n1183), .A3(n1487), .Z(N15154) );
  an02d0 U11809 ( .A1(n1298), .A2(n1243), .Z(n1488) );
  nd02d0 U11810 ( .A1(n1205), .A2(n1488), .ZN(n1491) );
  nd04d0 U11811 ( .A1(n1096), .A2(n1072), .A3(n1025), .A4(n981), .ZN(n1490) );
  aoi21d1 U11812 ( .B1(n1141), .B2(n1488), .A(n1492), .ZN(n1489) );
  aoi211d1 U11813 ( .C1(n1491), .C2(n1490), .A(n1361), .B(n1489), .ZN(N15122)
         );
  an02d0 U11814 ( .A1(n1338), .A2(n1296), .Z(n1495) );
  an03d0 U11815 ( .A1(n1070), .A2(n1021), .A3(n1093), .Z(n1493) );
  nd04d0 U11816 ( .A1(n1495), .A2(n1142), .A3(n1254), .A4(n1493), .ZN(n1494)
         );
  oaim31d1 U11817 ( .B1(n1231), .B2(n1495), .B3(n1188), .A(n1494), .ZN(N15106)
         );
  an02d0 U11818 ( .A1(n1298), .A2(n1243), .Z(n1496) );
  nd02d0 U11819 ( .A1(n1205), .A2(n1496), .ZN(n1499) );
  oai211d1 U11820 ( .C1(n961), .C2(n999), .A(n1066), .B(n1096), .ZN(n1498) );
  aoi21d1 U11821 ( .B1(n1142), .B2(n1496), .A(n1500), .ZN(n1497) );
  aoi211d1 U11822 ( .C1(n1499), .C2(n1498), .A(n1361), .B(n1497), .ZN(N15090)
         );
  aor31d1 U11823 ( .B1(n1110), .B2(n1064), .B3(n1136), .A(n1194), .Z(n1501) );
  an04d0 U11824 ( .A1(n1342), .A2(n1300), .A3(n1246), .A4(n1501), .Z(N15074)
         );
  an02d0 U11825 ( .A1(n1298), .A2(n1243), .Z(n1502) );
  an02d0 U11826 ( .A1(n1201), .A2(n1502), .Z(n1503) );
  aoi21d1 U11827 ( .B1(n1142), .B2(n1502), .A(n1503), .ZN(n1505) );
  aoi321d1 U11828 ( .C1(n972), .C2(n1091), .C3(n1018), .B1(n1109), .B2(n1054), 
        .A(n1503), .ZN(n1504) );
  nr13d1 U11829 ( .A1(n1343), .A2(n1505), .A3(n1504), .ZN(N15058) );
  oai211d1 U11830 ( .C1(n998), .C2(n1044), .A(n1111), .B(n1139), .ZN(n1508) );
  nd02d0 U11831 ( .A1(n1345), .A2(n1305), .ZN(n1507) );
  nd13d1 U11832 ( .A1(n1507), .A2(n1238), .A3(n1178), .ZN(n1506) );
  oai31d1 U11833 ( .B1(n1508), .B2(n1507), .B3(n1267), .A(n1506), .ZN(N15042)
         );
  an02d0 U11834 ( .A1(n1297), .A2(n1243), .Z(n1510) );
  an02d0 U11835 ( .A1(n1200), .A2(n1510), .Z(n1509) );
  aoi21d1 U11836 ( .B1(n1100), .B2(n1049), .A(n1509), .ZN(n1513) );
  oai21d1 U11837 ( .B1(n972), .B2(n1011), .A(n1103), .ZN(n1512) );
  aoi21d1 U11838 ( .B1(n1142), .B2(n1510), .A(n1509), .ZN(n1511) );
  aoi211d1 U11839 ( .C1(n1513), .C2(n1512), .A(n1361), .B(n1511), .ZN(N15026)
         );
  aon211d1 U11840 ( .C1(n1139), .C2(n1089), .B(n1204), .A(n1233), .ZN(n1514)
         );
  nr23d1 U11841 ( .A1(n1334), .A2(n1294), .A3(n1514), .ZN(N15010) );
  an02d0 U11842 ( .A1(n1297), .A2(n1243), .Z(n1515) );
  an02d0 U11843 ( .A1(n1200), .A2(n1515), .Z(n1516) );
  aoi21d1 U11844 ( .B1(n1142), .B2(n1515), .A(n1516), .ZN(n1518) );
  aoi311d1 U11845 ( .C1(n1001), .C2(n962), .C3(n1043), .A(n1093), .B(n1516), 
        .ZN(n1517) );
  nr13d1 U11846 ( .A1(n1343), .A2(n1518), .A3(n1517), .ZN(N14994) );
  aoi31d1 U11847 ( .B1(n1068), .B2(n1015), .B3(n1148), .A(n1187), .ZN(n1519)
         );
  oaim21d1 U11848 ( .B1(n1115), .B2(n1138), .A(n1519), .ZN(n1520) );
  an02d0 U11849 ( .A1(n1298), .A2(n1243), .Z(n1521) );
  nd02d0 U11850 ( .A1(n1205), .A2(n1521), .ZN(n1524) );
  oai21d1 U11851 ( .B1(n972), .B2(n1011), .A(n1061), .ZN(n1523) );
  aoi21d1 U11852 ( .B1(n1143), .B2(n1521), .A(n1525), .ZN(n1522) );
  aoi311d1 U11853 ( .C1(n1524), .C2(n1128), .C3(n1523), .A(n1360), .B(n1522), 
        .ZN(N14962) );
  an04d0 U11854 ( .A1(n1342), .A2(n1300), .A3(n1246), .A4(n1999), .Z(N14946)
         );
  an02d0 U11855 ( .A1(n1298), .A2(n1243), .Z(n1527) );
  nd02d0 U11856 ( .A1(n1205), .A2(n1527), .ZN(n1526) );
  oaim21d1 U11857 ( .B1(n1020), .B2(n983), .A(n1526), .ZN(n1529) );
  oaim21d1 U11858 ( .B1(n1156), .B2(n1527), .A(n1526), .ZN(n1528) );
  ora311d1 U11859 ( .C1(n1113), .C2(n1045), .C3(n1529), .A(n1528), .B(n1334), 
        .Z(N14930) );
  oan211d1 U11860 ( .C1(n1007), .C2(n1049), .B(n1137), .A(n1189), .ZN(n1530)
         );
  oaim21d1 U11861 ( .B1(n1115), .B2(n1136), .A(n1530), .ZN(n1531) );
  nr02d0 U11862 ( .A1(n1026), .A2(n978), .ZN(n1533) );
  nr03d0 U11863 ( .A1(n1070), .A2(n1206), .A3(n1101), .ZN(n1532) );
  aoim22d1 U11864 ( .A1(n1533), .A2(n1532), .B1(n1198), .B2(n1152), .Z(n1534)
         );
  oai21d1 U11865 ( .B1(n1145), .B2(n1189), .A(n1234), .ZN(n1535) );
  nr23d1 U11866 ( .A1(n1324), .A2(n1304), .A3(n1535), .ZN(N14882) );
  an02d0 U11867 ( .A1(n1019), .A2(n978), .Z(n1536) );
  aor311d1 U11868 ( .C1(n1112), .C2(n1064), .C3(n1536), .A(n1205), .B(n1134), 
        .Z(n1537) );
  an04d0 U11869 ( .A1(n1341), .A2(n1300), .A3(n1247), .A4(n1537), .Z(N14866)
         );
  aor311d1 U11870 ( .C1(n1068), .C2(n1015), .C3(n1092), .A(n1200), .B(n1134), 
        .Z(n1538) );
  an04d0 U11871 ( .A1(n1342), .A2(n1299), .A3(n1246), .A4(n1538), .Z(N14850)
         );
  or02d0 U11872 ( .A1(n983), .A2(n1021), .Z(n1539) );
  aor311d1 U11873 ( .C1(n1068), .C2(n1539), .C3(n1092), .A(n1189), .B(n1135), 
        .Z(n1540) );
  an04d0 U11874 ( .A1(n1342), .A2(n1299), .A3(n1246), .A4(n1540), .Z(N14834)
         );
  aor211d1 U11875 ( .C1(n1111), .C2(n1050), .A(n1179), .B(n1156), .Z(n1541) );
  nd03d0 U11876 ( .A1(n982), .A2(n1096), .A3(n1028), .ZN(n1543) );
  nr02d0 U11877 ( .A1(n1207), .A2(n1160), .ZN(n1542) );
  oaim211d1 U11878 ( .C1(n1113), .C2(n1067), .A(n1543), .B(n1542), .ZN(n1544)
         );
  an04d0 U11879 ( .A1(n1342), .A2(n1299), .A3(n1246), .A4(n1544), .Z(N14802)
         );
  or02d0 U11880 ( .A1(n1028), .A2(n1082), .Z(n1545) );
  aor211d1 U11881 ( .C1(n1111), .C2(n1545), .A(n1179), .B(n1136), .Z(n1546) );
  oai21d1 U11882 ( .B1(n971), .B2(n1010), .A(n1103), .ZN(n1548) );
  nr02d0 U11883 ( .A1(n1189), .A2(n1160), .ZN(n1547) );
  oaim211d1 U11884 ( .C1(n1113), .C2(n1067), .A(n1548), .B(n1547), .ZN(n1549)
         );
  an04d0 U11885 ( .A1(n1341), .A2(n1299), .A3(n1247), .A4(n1549), .Z(N14770)
         );
  oai21d1 U11886 ( .B1(n1102), .B2(n1139), .A(n1228), .ZN(n1550) );
  oaim21d1 U11887 ( .B1(n1201), .B2(n1236), .A(n1550), .ZN(n1551) );
  an03d0 U11888 ( .A1(n1308), .A2(n1551), .A3(n1340), .Z(N14754) );
  aor31d1 U11889 ( .B1(n1018), .B2(n977), .B3(n1052), .A(n1106), .Z(n1553) );
  an02d0 U11890 ( .A1(n1338), .A2(n1295), .Z(n1552) );
  ora311d1 U11891 ( .C1(n1208), .C2(n1143), .C3(n1553), .A(n1244), .B(n1552), 
        .Z(N14738) );
  aoi211d1 U11892 ( .C1(n1062), .C2(n1008), .A(n1146), .B(n1089), .ZN(n1556)
         );
  nd02d0 U11893 ( .A1(n1345), .A2(n1304), .ZN(n1555) );
  nd13d1 U11894 ( .A1(n1555), .A2(n1238), .A3(n1207), .ZN(n1554) );
  oai31d1 U11895 ( .B1(n1259), .B2(n1556), .B3(n1555), .A(n1554), .ZN(N14722)
         );
  oan211d1 U11896 ( .C1(n966), .C2(n1003), .B(n1057), .A(n1097), .ZN(n1558) );
  nr02d0 U11897 ( .A1(n1180), .A2(n1160), .ZN(n1557) );
  nd02d0 U11898 ( .A1(n1558), .A2(n1557), .ZN(n1559) );
  an04d0 U11899 ( .A1(n1341), .A2(n1299), .A3(n1247), .A4(n1559), .Z(N14706)
         );
  or04d0 U11900 ( .A1(n1117), .A2(n1056), .A3(n1194), .A4(n1147), .Z(n1560) );
  an04d0 U11901 ( .A1(n1342), .A2(n1299), .A3(n1247), .A4(n1560), .Z(N14690)
         );
  aoi21d1 U11902 ( .B1(n1012), .B2(n964), .A(n1063), .ZN(n1562) );
  nr03d0 U11903 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n1561) );
  nd02d0 U11904 ( .A1(n1562), .A2(n1561), .ZN(n1563) );
  nr04d0 U11905 ( .A1(n1158), .A2(n1118), .A3(n1041), .A4(n1023), .ZN(n1566)
         );
  nd02d0 U11906 ( .A1(n1345), .A2(n1304), .ZN(n1565) );
  nd13d1 U11907 ( .A1(n1565), .A2(n1238), .A3(n1190), .ZN(n1564) );
  oai31d1 U11908 ( .B1(n1265), .B2(n1566), .B3(n1565), .A(n1564), .ZN(N14658)
         );
  nr03d0 U11909 ( .A1(n979), .A2(n1071), .A3(n1027), .ZN(n1568) );
  nr03d0 U11910 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n1567) );
  nd02d0 U11911 ( .A1(n1568), .A2(n1567), .ZN(n1569) );
  an03d0 U11912 ( .A1(n1308), .A2(n1248), .A3(n1339), .Z(N14626) );
  nd02d0 U11913 ( .A1(n1309), .A2(n1249), .ZN(n1572) );
  nd04d0 U11914 ( .A1(n1102), .A2(n1072), .A3(n1025), .A4(n980), .ZN(n1571) );
  aoi31d1 U11915 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n1527), .ZN(n1570)
         );
  aoi211d1 U11916 ( .C1(n1572), .C2(n1571), .A(n1361), .B(n1570), .ZN(N14610)
         );
  nd04d0 U11917 ( .A1(n1162), .A2(n1092), .A3(n1084), .A4(n1023), .ZN(n1573)
         );
  aoim22d1 U11918 ( .A1(n1573), .A2(n1259), .B1(n1198), .B2(n1238), .Z(n1574)
         );
  an03d0 U11919 ( .A1(n1345), .A2(n1301), .A3(n1574), .Z(N14594) );
  nd02d0 U11920 ( .A1(n1309), .A2(n1249), .ZN(n1577) );
  oai211d1 U11921 ( .C1(n961), .C2(n1023), .A(n1065), .B(n1097), .ZN(n1576) );
  aoi31d1 U11922 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n2238), .ZN(n1575)
         );
  aoi211d1 U11923 ( .C1(n1577), .C2(n1576), .A(n1361), .B(n1575), .ZN(N14578)
         );
  an03d0 U11924 ( .A1(n1118), .A2(n1076), .A3(n1156), .Z(n1578) );
  nd04d0 U11925 ( .A1(n1299), .A2(n1208), .A3(n1348), .A4(n1578), .ZN(n1579)
         );
  oaim31d1 U11926 ( .B1(n1334), .B2(n1288), .B3(n1237), .A(n1579), .ZN(N14562)
         );
  an02d0 U11927 ( .A1(n1244), .A2(n1296), .Z(n1580) );
  aoi31d1 U11928 ( .B1(n1196), .B2(n1151), .B3(n1285), .A(n1580), .ZN(n1582)
         );
  aoi321d1 U11929 ( .C1(n971), .C2(n1091), .C3(n1025), .B1(n1109), .B2(n1055), 
        .A(n1580), .ZN(n1581) );
  nr13d1 U11930 ( .A1(n1343), .A2(n1582), .A3(n1581), .ZN(N14546) );
  oai211d1 U11931 ( .C1(n1006), .C2(n1044), .A(n1110), .B(n1140), .ZN(n1583)
         );
  aoim22d1 U11932 ( .A1(n1583), .A2(n1266), .B1(n1197), .B2(n1238), .Z(n1584)
         );
  an03d0 U11933 ( .A1(n1345), .A2(n1301), .A3(n1584), .Z(N14530) );
  oai21d1 U11934 ( .B1(n971), .B2(n1011), .A(n1104), .ZN(n1588) );
  nd02d0 U11935 ( .A1(n1111), .A2(n1084), .ZN(n1587) );
  nd02d0 U11936 ( .A1(n1253), .A2(n1304), .ZN(n1586) );
  aoi31d1 U11937 ( .B1(n1196), .B2(n1151), .B3(n1285), .A(n1580), .ZN(n1585)
         );
  aoi311d1 U11938 ( .C1(n1588), .C2(n1587), .C3(n1586), .A(n1360), .B(n1585), 
        .ZN(N14514) );
  aor31d1 U11939 ( .B1(n1154), .B2(n1110), .B3(n1187), .A(n1235), .Z(n1589) );
  an03d0 U11940 ( .A1(n1308), .A2(n1589), .A3(n1340), .Z(N14498) );
  an02d0 U11941 ( .A1(n1244), .A2(n1296), .Z(n1590) );
  aoi31d1 U11942 ( .B1(n1196), .B2(n1151), .B3(n1286), .A(n1590), .ZN(n1592)
         );
  aoi311d1 U11943 ( .C1(n1027), .C2(n962), .C3(n1043), .A(n1590), .B(n1091), 
        .ZN(n1591) );
  nr13d1 U11944 ( .A1(n1343), .A2(n1592), .A3(n1591), .ZN(N14482) );
  nd02d0 U11945 ( .A1(n1345), .A2(n1304), .ZN(n1594) );
  aoi321d1 U11946 ( .C1(n1060), .C2(n1002), .C3(n1134), .B1(n1108), .B2(n1136), 
        .A(n1240), .ZN(n1593) );
  aoim211d1 U11947 ( .C1(n1188), .C2(n1227), .A(n1594), .B(n1593), .ZN(N14466)
         );
  oan211d1 U11948 ( .C1(n966), .C2(n1003), .B(n1056), .A(n1098), .ZN(n1597) );
  nd02d0 U11949 ( .A1(n1253), .A2(n1304), .ZN(n1596) );
  aoi31d1 U11950 ( .B1(n1196), .B2(n1151), .B3(n1286), .A(n1590), .ZN(n1595)
         );
  aoi211d1 U11951 ( .C1(n1597), .C2(n1596), .A(n1368), .B(n1595), .ZN(N14450)
         );
  ora211d1 U11952 ( .C1(n1046), .C2(n1101), .A(n1157), .B(n1199), .Z(n1598) );
  ora211d1 U11953 ( .C1(n1243), .C2(n1598), .A(n1301), .B(n1337), .Z(N14434)
         );
  nd02d0 U11954 ( .A1(n1309), .A2(n1249), .ZN(n1599) );
  oaim21d1 U11955 ( .B1(n1020), .B2(N6867), .A(n1599), .ZN(n1601) );
  oaim31d1 U11956 ( .B1(n1139), .B2(n1288), .B3(n1177), .A(n1599), .ZN(n1600)
         );
  ora311d1 U11957 ( .C1(n1109), .C2(n1045), .C3(n1601), .A(n1600), .B(n1335), 
        .Z(N14418) );
  oan211d1 U11958 ( .C1(n1007), .C2(n1048), .B(n1139), .A(n1232), .ZN(n1603)
         );
  nd02d0 U11959 ( .A1(n1094), .A2(n1159), .ZN(n1602) );
  aoim22d1 U11960 ( .A1(n1603), .A2(n1602), .B1(n1198), .B2(n1238), .Z(n1604)
         );
  an03d0 U11961 ( .A1(n1345), .A2(n1301), .A3(n1604), .Z(N14402) );
  nd02d0 U11962 ( .A1(n1309), .A2(n1248), .ZN(n1607) );
  nr03d0 U11963 ( .A1(n1021), .A2(n1119), .A3(n1037), .ZN(n1606) );
  aoi31d1 U11964 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n2123), .ZN(n1605)
         );
  aoi311d1 U11965 ( .C1(n1607), .C2(n992), .C3(n1606), .A(n1359), .B(n1605), 
        .ZN(N14386) );
  aon211d1 U11966 ( .C1(n1203), .C2(n1135), .B(n1225), .A(n1284), .ZN(n1608)
         );
  nr02d0 U11967 ( .A1(n1368), .A2(n1608), .ZN(N14370) );
  nd03d0 U11968 ( .A1(n1207), .A2(num_images[4]), .A3(n1286), .ZN(n1609) );
  oaim21d1 U11969 ( .B1(n1245), .B2(n1287), .A(n1609), .ZN(n1610) );
  nd04d0 U11970 ( .A1(n1119), .A2(n1072), .A3(n1024), .A4(n981), .ZN(n1612) );
  aoi21d1 U11971 ( .B1(n1279), .B2(n1187), .A(n1610), .ZN(n1611) );
  aoi211d1 U11972 ( .C1(n1613), .C2(n1612), .A(n1369), .B(n1611), .ZN(N14354)
         );
  nd02d0 U11973 ( .A1(n1345), .A2(n1304), .ZN(n1615) );
  aoi311d1 U11974 ( .C1(n1046), .C2(n1022), .C3(n1111), .A(n1229), .B(n1149), 
        .ZN(n1614) );
  aoim211d1 U11975 ( .C1(n1177), .C2(n1227), .A(n1615), .B(n1614), .ZN(N14338)
         );
  nd03d0 U11976 ( .A1(n1207), .A2(n1160), .A3(n1284), .ZN(n1616) );
  oaim21d1 U11977 ( .B1(n1245), .B2(n1276), .A(n1616), .ZN(n1617) );
  oai211d1 U11978 ( .C1(n960), .C2(n1025), .A(n1065), .B(n1097), .ZN(n1619) );
  aoi21d1 U11979 ( .B1(n1279), .B2(n1185), .A(n1617), .ZN(n1618) );
  aoi211d1 U11980 ( .C1(n1620), .C2(n1619), .A(n1356), .B(n1618), .ZN(N14322)
         );
  aoi321d1 U11981 ( .C1(n1101), .C2(n1047), .C3(n1177), .B1(n1148), .B2(n1188), 
        .A(n1241), .ZN(n1621) );
  nr23d1 U11982 ( .A1(n1283), .A2(n1350), .A3(n1621), .ZN(N14306) );
  nd03d0 U11983 ( .A1(n1207), .A2(n1140), .A3(n1274), .ZN(n1622) );
  oaim21d1 U11984 ( .B1(n1244), .B2(n1287), .A(n1622), .ZN(n1624) );
  aoi321d1 U11985 ( .C1(n971), .C2(n1091), .C3(n1023), .B1(n1107), .B2(n1054), 
        .A(n1624), .ZN(n1623) );
  aon211d1 U11986 ( .C1(n1180), .C2(n1283), .B(n1624), .A(n1626), .ZN(n1625)
         );
  nr02d0 U11987 ( .A1(n1625), .A2(n1371), .ZN(N14290) );
  nr02d0 U11988 ( .A1(n1255), .A2(n1160), .ZN(n1628) );
  oai21d1 U11989 ( .B1(n1012), .B2(n1058), .A(n1104), .ZN(n1627) );
  aoim22d1 U11990 ( .A1(n1628), .A2(n1627), .B1(n1197), .B2(n1237), .Z(n1629)
         );
  an03d0 U11991 ( .A1(n1345), .A2(n1301), .A3(n1629), .Z(N14274) );
  nd03d0 U11992 ( .A1(n1207), .A2(n1155), .A3(n1270), .ZN(n1630) );
  oaim21d1 U11993 ( .B1(n1245), .B2(n1287), .A(n1630), .ZN(n1633) );
  oai21d1 U11994 ( .B1(n971), .B2(n1009), .A(n1104), .ZN(n1631) );
  oaim2m11d1 U11995 ( .C1(n1114), .C2(n1064), .B(n1633), .A(n1631), .ZN(n1632)
         );
  aon211d1 U11996 ( .C1(n1180), .C2(n1304), .B(n1633), .A(n1632), .ZN(n1634)
         );
  nr02d0 U11997 ( .A1(n1634), .A2(n1367), .ZN(N14258) );
  oan211d1 U11998 ( .C1(n1092), .C2(n1132), .B(n1188), .A(n1232), .ZN(n1635)
         );
  nr23d1 U11999 ( .A1(n1302), .A2(n1350), .A3(n1635), .ZN(N14242) );
  nd03d0 U12000 ( .A1(n1207), .A2(n1156), .A3(n1283), .ZN(n1636) );
  oaim21d1 U12001 ( .B1(n1245), .B2(n1287), .A(n1636), .ZN(n1638) );
  aor311d1 U12002 ( .C1(n1017), .C2(n976), .C3(n1050), .A(n1638), .B(n1117), 
        .Z(n1637) );
  aon211d1 U12003 ( .C1(n1182), .C2(n1281), .B(n1638), .A(n1637), .ZN(n1639)
         );
  nr02d0 U12004 ( .A1(n1639), .A2(n1366), .ZN(N14226) );
  aoi21d1 U12005 ( .B1(n1059), .B2(n1005), .A(n1109), .ZN(n1641) );
  nr02d0 U12006 ( .A1(n1254), .A2(n1160), .ZN(n1640) );
  aoim22d1 U12007 ( .A1(n1641), .A2(n1640), .B1(n1197), .B2(n1238), .Z(n1642)
         );
  an03d0 U12008 ( .A1(n1345), .A2(n1301), .A3(n1642), .Z(N14210) );
  oan211d1 U12009 ( .C1(n966), .C2(n1004), .B(n1056), .A(n1099), .ZN(n1646) );
  nd03d0 U12010 ( .A1(n1207), .A2(n1135), .A3(n1287), .ZN(n1643) );
  oaim21d1 U12011 ( .B1(n1245), .B2(n1288), .A(n1643), .ZN(n1644) );
  aoi21d1 U12012 ( .B1(n1279), .B2(n1185), .A(n1644), .ZN(n1645) );
  aoi211d1 U12013 ( .C1(n1646), .C2(n1647), .A(n1368), .B(n1645), .ZN(N14194)
         );
  oan211d1 U12014 ( .C1(n1052), .C2(num_images[3]), .B(n1188), .A(n1232), .ZN(
        n1648) );
  oaim21d1 U12015 ( .B1(n1156), .B2(n1193), .A(n1648), .ZN(n1649) );
  an03d0 U12016 ( .A1(n1307), .A2(n1649), .A3(n1339), .Z(N14178) );
  an03d0 U12017 ( .A1(n1204), .A2(n1157), .A3(n1300), .Z(n1650) );
  aoi21d1 U12018 ( .B1(n1233), .B2(n1273), .A(n1650), .ZN(n1651) );
  oaim21d1 U12019 ( .B1(n1020), .B2(n957), .A(n1651), .ZN(n1653) );
  oaim21d1 U12020 ( .B1(n1201), .B2(n1288), .A(n1651), .ZN(n1652) );
  ora311d1 U12021 ( .C1(n1093), .C2(n1045), .C3(n1653), .A(n1652), .B(n1334), 
        .Z(N14162) );
  nr02d0 U12022 ( .A1(n1085), .A2(n1021), .ZN(n1655) );
  nr03d0 U12023 ( .A1(n1118), .A2(n1253), .A3(n1163), .ZN(n1654) );
  aoim22d1 U12024 ( .A1(n1655), .A2(n1654), .B1(n1198), .B2(n1237), .Z(n1656)
         );
  an03d0 U12025 ( .A1(n1345), .A2(n1300), .A3(n1656), .Z(N14146) );
  nd03d0 U12026 ( .A1(n1207), .A2(n1162), .A3(n1275), .ZN(n1657) );
  oaim21d1 U12027 ( .B1(n1246), .B2(n1288), .A(n1657), .ZN(n1660) );
  or03d0 U12028 ( .A1(n1089), .A2(n1081), .A3(n1020), .Z(n1659) );
  aor21d1 U12029 ( .B1(n1200), .B2(n1279), .A(n1660), .Z(n1658) );
  ora311d1 U12030 ( .C1(n963), .C2(n1660), .C3(n1659), .A(n1658), .B(n1335), 
        .Z(N14130) );
  ora211d1 U12031 ( .C1(n1184), .C2(n1234), .A(n1301), .B(n1337), .Z(N14114)
         );
  aoi22d1 U12032 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1177), .ZN(n1663)
         );
  nd04d0 U12033 ( .A1(n1120), .A2(n1072), .A3(n1024), .A4(n981), .ZN(n1662) );
  aoi21d1 U12034 ( .B1(n1144), .B2(n1273), .A(n1677), .ZN(n1661) );
  aoi211d1 U12035 ( .C1(n1663), .C2(n1662), .A(n1370), .B(n1661), .ZN(N14098)
         );
  an04d0 U12036 ( .A1(n1159), .A2(n1115), .A3(n1054), .A4(n1019), .Z(n1664) );
  ora311d1 U12037 ( .C1(n1224), .C2(n1178), .C3(n1664), .A(n1297), .B(n1335), 
        .Z(N14082) );
  aoi22d1 U12038 ( .A1(n1226), .A2(n1272), .B1(n1284), .B2(n1177), .ZN(n1667)
         );
  oai211d1 U12039 ( .C1(n960), .C2(n999), .A(n1066), .B(n1097), .ZN(n1666) );
  aoi21d1 U12040 ( .B1(n1143), .B2(n1273), .A(n2328), .ZN(n1665) );
  aoi211d1 U12041 ( .C1(n1667), .C2(n1666), .A(n1366), .B(n1665), .ZN(N14066)
         );
  aor311d1 U12042 ( .C1(n1112), .C2(n1064), .C3(n1155), .A(n1223), .B(n1178), 
        .Z(n1668) );
  an03d0 U12043 ( .A1(n1308), .A2(n1668), .A3(n1339), .Z(N14050) );
  aor22d1 U12044 ( .A1(n1238), .A2(n1282), .B1(n1292), .B2(n1179), .Z(n1669)
         );
  aoi321d1 U12045 ( .C1(n970), .C2(n1087), .C3(n1000), .B1(n1108), .B2(n1054), 
        .A(n1669), .ZN(n1671) );
  aoi21d1 U12046 ( .B1(n1144), .B2(n1273), .A(n1669), .ZN(n1670) );
  nr13d1 U12047 ( .A1(n1343), .A2(n1671), .A3(n1670), .ZN(N14034) );
  ora211d1 U12048 ( .C1(n1002), .C2(n1060), .A(n1116), .B(n1155), .Z(n1672) );
  ora311d1 U12049 ( .C1(n1224), .C2(n1178), .C3(n1672), .A(n1296), .B(n1335), 
        .Z(N14018) );
  oai21d1 U12050 ( .B1(n970), .B2(n1009), .A(n1105), .ZN(n1676) );
  nd02d0 U12051 ( .A1(n1110), .A2(n1085), .ZN(n1675) );
  aoi22d1 U12052 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1177), .ZN(n1674)
         );
  aoi21d1 U12053 ( .B1(n1144), .B2(n1273), .A(n1677), .ZN(n1673) );
  aoi311d1 U12054 ( .C1(n1676), .C2(n1675), .C3(n1674), .A(n1360), .B(n1673), 
        .ZN(N14002) );
  aor211d1 U12055 ( .C1(n1153), .C2(n1092), .A(n1237), .B(n1181), .Z(n1678) );
  an03d0 U12056 ( .A1(n1308), .A2(n1340), .A3(n1678), .Z(N13986) );
  aor22d1 U12057 ( .A1(n1238), .A2(n1282), .B1(n1292), .B2(n1179), .Z(n1679)
         );
  aoi311d1 U12058 ( .C1(n1001), .C2(n962), .C3(n1043), .A(n1679), .B(n1118), 
        .ZN(n1681) );
  aoi21d1 U12059 ( .B1(n1143), .B2(n1273), .A(n1679), .ZN(n1680) );
  nr13d1 U12060 ( .A1(n1343), .A2(n1681), .A3(n1680), .ZN(N13970) );
  nd03d0 U12061 ( .A1(n1071), .A2(n1028), .A3(n1163), .ZN(n1682) );
  oaim21d1 U12062 ( .B1(n1115), .B2(n1148), .A(n1682), .ZN(n1683) );
  ora311d1 U12063 ( .C1(n1224), .C2(n1179), .C3(n1683), .A(n1297), .B(n1335), 
        .Z(N13954) );
  oan211d1 U12064 ( .C1(n965), .C2(n1004), .B(n1056), .A(n1100), .ZN(n1686) );
  aoi22d1 U12065 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1177), .ZN(n1685)
         );
  aoi21d1 U12066 ( .B1(n1143), .B2(n1273), .A(n1677), .ZN(n1684) );
  aoi211d1 U12067 ( .C1(n1686), .C2(n1685), .A(n1360), .B(n1684), .ZN(N13938)
         );
  oai21d1 U12068 ( .B1(n1060), .B2(n1097), .A(n1146), .ZN(n1687) );
  ora311d1 U12069 ( .C1(n1224), .C2(n1178), .C3(n1688), .A(n1297), .B(n1334), 
        .Z(N13922) );
  aoi22d1 U12070 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1177), .ZN(n1689)
         );
  oaim21d1 U12071 ( .B1(n1020), .B2(n975), .A(n1689), .ZN(n1691) );
  oaim21d1 U12072 ( .B1(n1156), .B2(n1287), .A(n1689), .ZN(n1690) );
  ora311d1 U12073 ( .C1(n1112), .C2(n1044), .C3(n1691), .A(n1690), .B(n1336), 
        .Z(N13906) );
  oai21d1 U12074 ( .B1(n1013), .B2(n1058), .A(n1146), .ZN(n1692) );
  oaim21d1 U12075 ( .B1(n1115), .B2(n1147), .A(n1692), .ZN(n1693) );
  ora311d1 U12076 ( .C1(n1224), .C2(n1178), .C3(n1693), .A(n1297), .B(n1335), 
        .Z(N13890) );
  aoi22d1 U12077 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1177), .ZN(n1696)
         );
  nr03d0 U12078 ( .A1(n1021), .A2(n1119), .A3(n1083), .ZN(n1695) );
  aoi21d1 U12079 ( .B1(n1144), .B2(n1297), .A(n1677), .ZN(n1694) );
  aoi311d1 U12080 ( .C1(n1696), .C2(n992), .C3(n1695), .A(n1359), .B(n1694), 
        .ZN(N13874) );
  oai21d1 U12081 ( .B1(n1145), .B2(n1188), .A(n1281), .ZN(n1697) );
  aon211d1 U12082 ( .C1(n1225), .C2(n1275), .B(n1699), .A(n1331), .ZN(n1698)
         );
  nd04d0 U12083 ( .A1(n1103), .A2(n1086), .A3(n1024), .A4(n981), .ZN(n1700) );
  nd12d0 U12084 ( .A1(n1163), .A2(n1700), .ZN(n1701) );
  aor31d1 U12085 ( .B1(n1069), .B2(n1016), .B3(n1092), .A(n1147), .Z(n1702) );
  ora311d1 U12086 ( .C1(n1249), .C2(n1179), .C3(n1702), .A(n1296), .B(n1335), 
        .Z(N13826) );
  oai211d1 U12087 ( .C1(n960), .C2(n999), .A(n1066), .B(n1097), .ZN(n1703) );
  nd12d0 U12088 ( .A1(n1162), .A2(n1703), .ZN(n1704) );
  ora311d1 U12089 ( .C1(n1224), .C2(n1179), .C3(n1704), .A(n1297), .B(n1335), 
        .Z(N13810) );
  aor21d1 U12090 ( .B1(n1112), .B2(n1060), .A(n1145), .Z(n1705) );
  ora311d1 U12091 ( .C1(n1224), .C2(n1178), .C3(n1705), .A(n1297), .B(n1336), 
        .Z(N13794) );
  nd03d0 U12092 ( .A1(n982), .A2(n1113), .A3(n1028), .ZN(n1707) );
  nr03d0 U12093 ( .A1(n1160), .A2(n1253), .A3(n1175), .ZN(n1706) );
  oaim211d1 U12094 ( .C1(n1113), .C2(n1067), .A(n1707), .B(n1706), .ZN(n1708)
         );
  an03d0 U12095 ( .A1(n1308), .A2(n1708), .A3(n1339), .Z(N13778) );
  ora311d1 U12096 ( .C1(n1224), .C2(n1178), .C3(n1865), .A(n1296), .B(n1336), 
        .Z(N13762) );
  oai21d1 U12097 ( .B1(n970), .B2(n1010), .A(n1104), .ZN(n1710) );
  nr03d0 U12098 ( .A1(n1140), .A2(n1224), .A3(num_images[5]), .ZN(n1709) );
  oaim211d1 U12099 ( .C1(n1113), .C2(n1067), .A(n1710), .B(n1709), .ZN(n1711)
         );
  an03d0 U12100 ( .A1(n1308), .A2(n1711), .A3(n1339), .Z(N13746) );
  or04d0 U12101 ( .A1(n1229), .A2(n1200), .A3(n1153), .A4(n1105), .Z(n1712) );
  an03d0 U12102 ( .A1(n1309), .A2(n1325), .A3(n1712), .Z(N13730) );
  or02d0 U12103 ( .A1(n1254), .A2(n1184), .Z(n1714) );
  aor31d1 U12104 ( .B1(n1018), .B2(n977), .B3(n1052), .A(n1106), .Z(n1713) );
  ora311d1 U12105 ( .C1(n1144), .C2(n1714), .C3(n1713), .A(n1296), .B(n1336), 
        .Z(N13714) );
  aoi21d1 U12106 ( .B1(n1059), .B2(n1006), .A(n1109), .ZN(n1716) );
  nr03d0 U12107 ( .A1(n1158), .A2(n1253), .A3(n1209), .ZN(n1715) );
  oaim211d1 U12108 ( .C1(n1716), .C2(n1715), .A(n1292), .B(n1339), .ZN(n1717)
         );
  oan211d1 U12109 ( .C1(n967), .C2(n1004), .B(n1055), .A(n1098), .ZN(n1719) );
  nr03d0 U12110 ( .A1(n1157), .A2(n1237), .A3(n1188), .ZN(n1718) );
  oaim211d1 U12111 ( .C1(n1719), .C2(n1718), .A(n1292), .B(n1350), .ZN(n1720)
         );
  or03d0 U12112 ( .A1(n1244), .A2(n1202), .A3(n1157), .Z(n1721) );
  ora311d1 U12113 ( .C1(n1118), .C2(n1044), .C3(n1721), .A(n1296), .B(n1335), 
        .Z(N13666) );
  aoi211d1 U12114 ( .C1(n1014), .C2(n967), .A(n1102), .B(n1045), .ZN(n1723) );
  nr03d0 U12115 ( .A1(n1160), .A2(n1253), .A3(num_images[5]), .ZN(n1722) );
  oaim211d1 U12116 ( .C1(n1723), .C2(n1722), .A(n1292), .B(n1334), .ZN(n1724)
         );
  nr03d0 U12117 ( .A1(n1022), .A2(n1119), .A3(n1081), .ZN(n1726) );
  nr03d0 U12118 ( .A1(n1161), .A2(n1223), .A3(n1187), .ZN(n1725) );
  oaim211d1 U12119 ( .C1(n1726), .C2(n1725), .A(n1292), .B(n1349), .ZN(n1727)
         );
  nr03d0 U12120 ( .A1(n979), .A2(n1071), .A3(n1027), .ZN(n1729) );
  nr04d0 U12121 ( .A1(n1227), .A2(n1204), .A3(n1162), .A4(n1106), .ZN(n1728)
         );
  oaim211d1 U12122 ( .C1(n1729), .C2(n1728), .A(n1293), .B(n1324), .ZN(n1730)
         );
  an02d0 U12123 ( .A1(n1339), .A2(n1295), .Z(N13602) );
  nd04d0 U12124 ( .A1(n1120), .A2(n1072), .A3(n1024), .A4(n979), .ZN(n1732) );
  aoi31d1 U12125 ( .B1(n1196), .B2(n1149), .B3(n1235), .A(n1289), .ZN(n1731)
         );
  aoi211d1 U12126 ( .C1(n1732), .C2(n1319), .A(n1353), .B(n1731), .ZN(N13586)
         );
  nd04d0 U12127 ( .A1(n1146), .A2(n1112), .A3(n1077), .A4(n1023), .ZN(n1735)
         );
  nd02d0 U12128 ( .A1(n1309), .A2(n1341), .ZN(n1734) );
  nd03d0 U12129 ( .A1(n1241), .A2(n1208), .A3(n1338), .ZN(n1733) );
  aoi22d1 U12130 ( .A1(n1735), .A2(n1322), .B1(n1734), .B2(n1733), .ZN(N13570)
         );
  oai211d1 U12131 ( .C1(n960), .C2(n999), .A(n1066), .B(n1097), .ZN(n1737) );
  aoi31d1 U12132 ( .B1(n1196), .B2(n1150), .B3(n1236), .A(n1289), .ZN(n1736)
         );
  aoi211d1 U12133 ( .C1(n1737), .C2(n1319), .A(n1360), .B(n1736), .ZN(N13554)
         );
  nd04d0 U12134 ( .A1(n1189), .A2(n1137), .A3(n1094), .A4(n1071), .ZN(n1738)
         );
  aoim22d1 U12135 ( .A1(n1738), .A2(n1318), .B1(n1240), .B2(n1292), .Z(n1739)
         );
  an02d0 U12136 ( .A1(n1739), .A2(n1337), .Z(N13538) );
  aoi31d1 U12137 ( .B1(n1197), .B2(n1149), .B3(n1236), .A(n1289), .ZN(n1741)
         );
  aoi321d1 U12138 ( .C1(n970), .C2(n1090), .C3(n1000), .B1(n1108), .B2(n1053), 
        .A(n1294), .ZN(n1740) );
  nr13d1 U12139 ( .A1(n1343), .A2(n1741), .A3(n1740), .ZN(N13522) );
  oai211d1 U12140 ( .C1(n998), .C2(n1044), .A(n1111), .B(n1139), .ZN(n1744) );
  nd02d0 U12141 ( .A1(n1292), .A2(n1341), .ZN(n1743) );
  nd03d0 U12142 ( .A1(n1235), .A2(n1208), .A3(n1336), .ZN(n1742) );
  aoi22d1 U12143 ( .A1(n1744), .A2(n1323), .B1(n1743), .B2(n1742), .ZN(N13506)
         );
  aoi21d1 U12144 ( .B1(n1100), .B2(n1050), .A(n1288), .ZN(n1747) );
  oai21d1 U12145 ( .B1(n969), .B2(n1010), .A(n1103), .ZN(n1746) );
  aoi31d1 U12146 ( .B1(n1197), .B2(n1150), .B3(n1236), .A(n1288), .ZN(n1745)
         );
  aoi211d1 U12147 ( .C1(n1747), .C2(n1746), .A(n1360), .B(n1745), .ZN(N13490)
         );
  an04d0 U12148 ( .A1(n1249), .A2(n1201), .A3(n1157), .A4(n1112), .Z(n1748) );
  oai21d1 U12149 ( .B1(n1279), .B2(n1748), .A(n1329), .ZN(n1749) );
  aoi31d1 U12150 ( .B1(n1197), .B2(n1150), .B3(n1236), .A(n1288), .ZN(n1751)
         );
  aoi311d1 U12151 ( .C1(n1001), .C2(n963), .C3(n1043), .A(n1274), .B(n1089), 
        .ZN(n1750) );
  nr13d1 U12152 ( .A1(n1343), .A2(n1751), .A3(n1750), .ZN(N13458) );
  nd03d0 U12153 ( .A1(n1236), .A2(n1209), .A3(n1333), .ZN(n1753) );
  aoi321d1 U12154 ( .C1(n1060), .C2(n1003), .C3(n1160), .B1(n1109), .B2(n1136), 
        .A(n1294), .ZN(n1752) );
  oan211d1 U12155 ( .C1(n1358), .C2(n1322), .B(n1753), .A(n1752), .ZN(N13442)
         );
  oai21d1 U12156 ( .B1(n969), .B2(n1010), .A(n1062), .ZN(n1754) );
  aor31d1 U12157 ( .B1(n1199), .B2(n1151), .B3(n1229), .A(n1283), .Z(n1755) );
  ora311d1 U12158 ( .C1(n1090), .C2(n1291), .C3(n1756), .A(n1338), .B(n1755), 
        .Z(N13426) );
  oai211d1 U12159 ( .C1(n1042), .C2(n1114), .A(n1153), .B(n1188), .ZN(n1757)
         );
  aoim22d1 U12160 ( .A1(n1757), .A2(n1318), .B1(n1240), .B2(n1292), .Z(n1758)
         );
  an02d0 U12161 ( .A1(n1758), .A2(n1337), .Z(N13410) );
  aor21d1 U12162 ( .B1(n1018), .B2(n969), .A(n1061), .Z(n1760) );
  aor31d1 U12163 ( .B1(n1199), .B2(n1151), .B3(n1229), .A(n1283), .Z(n1759) );
  ora311d1 U12164 ( .C1(n1114), .C2(n1272), .C3(n1760), .A(n1338), .B(n1759), 
        .Z(N13394) );
  nd03d0 U12165 ( .A1(n1246), .A2(n1208), .A3(N11556), .ZN(n1763) );
  oai21d1 U12166 ( .B1(n1012), .B2(n1058), .A(n1147), .ZN(n1761) );
  aoi211d1 U12167 ( .C1(n1106), .C2(n1138), .A(n1281), .B(n1764), .ZN(n1762)
         );
  oan211d1 U12168 ( .C1(n1359), .C2(n1319), .B(n1763), .A(n1762), .ZN(N13378)
         );
  or03d0 U12169 ( .A1(n1295), .A2(n1117), .A3(n1053), .Z(n1766) );
  aor31d1 U12170 ( .B1(n1199), .B2(n1151), .B3(n1228), .A(n1283), .Z(n1765) );
  ora311d1 U12171 ( .C1(n1002), .C2(n963), .C3(n1766), .A(n1765), .B(n1335), 
        .Z(N13362) );
  aor31d1 U12172 ( .B1(n1198), .B2(n1152), .B3(n1229), .A(n1284), .Z(n1767) );
  an02d0 U12173 ( .A1(n1339), .A2(n1767), .Z(N13346) );
  aoi31d1 U12174 ( .B1(n1197), .B2(n1150), .B3(n1236), .A(n1286), .ZN(n1770)
         );
  nd04d0 U12175 ( .A1(n1120), .A2(n1037), .A3(n1025), .A4(n980), .ZN(n1769) );
  aoi21d1 U12176 ( .B1(n1234), .B2(n1185), .A(n1765), .ZN(n1768) );
  aoi211d1 U12177 ( .C1(n1770), .C2(n1769), .A(n1360), .B(n1768), .ZN(N13330)
         );
  nd03d0 U12178 ( .A1(n1240), .A2(n1208), .A3(n1340), .ZN(n1772) );
  aoi311d1 U12179 ( .C1(n1046), .C2(n1021), .C3(n1117), .A(n1274), .B(n1134), 
        .ZN(n1771) );
  oan211d1 U12180 ( .C1(n1359), .C2(n1310), .B(n1772), .A(n1771), .ZN(N13314)
         );
  aoi31d1 U12181 ( .B1(n1196), .B2(n1151), .B3(n1235), .A(n1288), .ZN(n1775)
         );
  oai211d1 U12182 ( .C1(n960), .C2(n1015), .A(n1065), .B(n1096), .ZN(n1774) );
  aoi21d1 U12183 ( .B1(n1233), .B2(n1185), .A(n1767), .ZN(n1773) );
  aoi211d1 U12184 ( .C1(n1775), .C2(n1774), .A(n1360), .B(n1773), .ZN(N13298)
         );
  aoi321d1 U12185 ( .C1(n1101), .C2(n1047), .C3(n1177), .B1(n1148), .B2(n1188), 
        .A(n1294), .ZN(n1776) );
  aoim2m11d1 U12186 ( .C1(n1234), .C2(n1309), .B(n1325), .A(n1776), .ZN(N13282) );
  aor31d1 U12187 ( .B1(n1199), .B2(n1152), .B3(n1228), .A(n1284), .Z(n1778) );
  aoi321d1 U12188 ( .C1(n969), .C2(n1087), .C3(n1000), .B1(n1107), .B2(n1053), 
        .A(n1778), .ZN(n1777) );
  aon211d1 U12189 ( .C1(n1180), .C2(n1251), .B(n1778), .A(n1780), .ZN(n1779)
         );
  nr02d0 U12190 ( .A1(n1779), .A2(n1356), .ZN(N13266) );
  nd03d0 U12191 ( .A1(n1243), .A2(n1209), .A3(n1339), .ZN(n1783) );
  or02d0 U12192 ( .A1(n1163), .A2(n1303), .Z(n1781) );
  oan211d1 U12193 ( .C1(n1007), .C2(n1048), .B(n1094), .A(n1781), .ZN(n1782)
         );
  oan211d1 U12194 ( .C1(n1358), .C2(n1271), .B(n1783), .A(n1782), .ZN(N13250)
         );
  aor31d1 U12195 ( .B1(n1199), .B2(n1152), .B3(n1228), .A(n1284), .Z(n1786) );
  oai21d1 U12196 ( .B1(n969), .B2(n1010), .A(n1103), .ZN(n1784) );
  oaim2m11d1 U12197 ( .C1(n1114), .C2(n1064), .B(n1786), .A(n1784), .ZN(n1785)
         );
  aon211d1 U12198 ( .C1(n1180), .C2(n1223), .B(n1786), .A(n1785), .ZN(n1787)
         );
  nr02d0 U12199 ( .A1(n1787), .A2(n1371), .ZN(N13234) );
  ora211d1 U12200 ( .C1(n1090), .C2(n1145), .A(n1207), .B(n1241), .Z(n1788) );
  oai21d1 U12201 ( .B1(n1279), .B2(n1788), .A(n1329), .ZN(n1789) );
  aor31d1 U12202 ( .B1(n1199), .B2(n1152), .B3(n1228), .A(n1283), .Z(n1791) );
  aor311d1 U12203 ( .C1(n1017), .C2(n976), .C3(n1050), .A(n1791), .B(n1098), 
        .Z(n1790) );
  aon211d1 U12204 ( .C1(n1183), .C2(n1245), .B(n1791), .A(n1790), .ZN(n1792)
         );
  nr02d0 U12205 ( .A1(n1792), .A2(n1367), .ZN(N13202) );
  nd03d0 U12206 ( .A1(n1231), .A2(n1208), .A3(n1337), .ZN(n1795) );
  or02d0 U12207 ( .A1(n1163), .A2(n1303), .Z(n1793) );
  aoi211d1 U12208 ( .C1(n1062), .C2(n1008), .A(n1793), .B(n1106), .ZN(n1794)
         );
  oan211d1 U12209 ( .C1(n1358), .C2(n1320), .B(n1795), .A(n1794), .ZN(N13186)
         );
  oan211d1 U12210 ( .C1(n967), .C2(n1005), .B(n1056), .A(n1097), .ZN(n1798) );
  aoi31d1 U12211 ( .B1(n1197), .B2(n1150), .B3(n1235), .A(n1289), .ZN(n1797)
         );
  aoi21d1 U12212 ( .B1(n1234), .B2(n1184), .A(n1759), .ZN(n1796) );
  aoi211d1 U12213 ( .C1(n1798), .C2(n1797), .A(n1360), .B(n1796), .ZN(N13170)
         );
  oan211d1 U12214 ( .C1(n1051), .C2(num_images[3]), .B(n1188), .A(n1276), .ZN(
        n1799) );
  oaim21d1 U12215 ( .B1(n1156), .B2(n1193), .A(n1799), .ZN(n1800) );
  aoi31d1 U12216 ( .B1(n1197), .B2(n1150), .B3(n1235), .A(n1289), .ZN(n1801)
         );
  oaim21d1 U12217 ( .B1(n1020), .B2(n975), .A(n1801), .ZN(n1803) );
  oaim21d1 U12218 ( .B1(n1201), .B2(n1237), .A(n1801), .ZN(n1802) );
  ora311d1 U12219 ( .C1(n1096), .C2(n1045), .C3(n1803), .A(n1802), .B(n1335), 
        .Z(N13138) );
  nd03d0 U12220 ( .A1(n1247), .A2(n1208), .A3(n1341), .ZN(n1806) );
  or02d0 U12221 ( .A1(n1163), .A2(n1303), .Z(n1804) );
  nr04d0 U12222 ( .A1(n1117), .A2(n1804), .A3(n1075), .A4(n1022), .ZN(n1805)
         );
  oan211d1 U12223 ( .C1(n1358), .C2(n1319), .B(n1806), .A(n1805), .ZN(N13122)
         );
  aoi31d1 U12224 ( .B1(n1196), .B2(n1150), .B3(n1235), .A(n1289), .ZN(n1809)
         );
  nr03d0 U12225 ( .A1(n1118), .A2(n1071), .A3(n1028), .ZN(n1808) );
  aoi21d1 U12226 ( .B1(n1190), .B2(n1221), .A(n1786), .ZN(n1807) );
  aoi311d1 U12227 ( .C1(n993), .C2(n1809), .C3(n1808), .A(n1807), .B(n1357), 
        .ZN(N13106) );
  nd03d0 U12228 ( .A1(n1229), .A2(n1209), .A3(N11556), .ZN(n1810) );
  oaim21d1 U12229 ( .B1(n1300), .B2(n1331), .A(n1810), .ZN(N13090) );
  aoi21d1 U12230 ( .B1(n1234), .B2(n1184), .A(n1289), .ZN(n1813) );
  nd04d0 U12231 ( .A1(n1120), .A2(n1080), .A3(n1024), .A4(n980), .ZN(n1812) );
  aoi21d1 U12232 ( .B1(n1143), .B2(n1244), .A(n1820), .ZN(n1811) );
  aoi211d1 U12233 ( .C1(n1813), .C2(n1812), .A(n1360), .B(n1811), .ZN(N13074)
         );
  an04d0 U12234 ( .A1(n1159), .A2(n1115), .A3(n1039), .A4(n1019), .Z(n1815) );
  aoi22d1 U12235 ( .A1(n1325), .A2(n1224), .B1(n1285), .B2(n1350), .ZN(n1814)
         );
  aoim31d1 U12236 ( .B1(n1189), .B2(n1273), .B3(n1815), .A(n1814), .ZN(N13058)
         );
  aoi21d1 U12237 ( .B1(n1233), .B2(n1185), .A(n1288), .ZN(n1818) );
  oai211d1 U12238 ( .C1(n961), .C2(n1018), .A(n1065), .B(n1095), .ZN(n1817) );
  aoi21d1 U12239 ( .B1(n1144), .B2(num_images[6]), .A(n2492), .ZN(n1816) );
  aoi211d1 U12240 ( .C1(n1818), .C2(n1817), .A(n1355), .B(n1816), .ZN(N13042)
         );
  aoi311d1 U12241 ( .C1(n1101), .C2(n1044), .C3(n1156), .A(n1274), .B(n1184), 
        .ZN(n1819) );
  aoim2m11d1 U12242 ( .C1(n1234), .C2(n1290), .B(n1332), .A(n1819), .ZN(N13026) );
  aor21d1 U12243 ( .B1(n1241), .B2(n1191), .A(n1280), .Z(n1820) );
  aoi321d1 U12244 ( .C1(n969), .C2(n1090), .C3(n1024), .B1(n1107), .B2(n1053), 
        .A(n1820), .ZN(n1822) );
  aoi21d1 U12245 ( .B1(n1144), .B2(n1243), .A(n1820), .ZN(n1821) );
  nr13d1 U12246 ( .A1(n1343), .A2(n1822), .A3(n1821), .ZN(N13010) );
  ora211d1 U12247 ( .C1(n1002), .C2(n1060), .A(n1116), .B(n1155), .Z(n1824) );
  aoi22d1 U12248 ( .A1(n1335), .A2(n1235), .B1(n1284), .B2(n1349), .ZN(n1823)
         );
  aoim31d1 U12249 ( .B1(num_images[5]), .B2(n1308), .B3(n1824), .A(n1823), 
        .ZN(N12994) );
  oai21d1 U12250 ( .B1(n968), .B2(n1009), .A(n1104), .ZN(n1828) );
  nd02d0 U12251 ( .A1(n1108), .A2(n1040), .ZN(n1827) );
  aoi21d1 U12252 ( .B1(n1233), .B2(n1184), .A(n1288), .ZN(n1826) );
  aoi21d1 U12253 ( .B1(n1144), .B2(n1246), .A(n1829), .ZN(n1825) );
  aoi311d1 U12254 ( .C1(n1828), .C2(n1827), .C3(n1826), .A(n1359), .B(n1825), 
        .ZN(N12978) );
  an03d0 U12255 ( .A1(n1100), .A2(n1248), .A3(n1157), .Z(n1830) );
  aon211d1 U12256 ( .C1(n1225), .C2(n1179), .B(n1830), .A(n1331), .ZN(n1831)
         );
  oaim21d1 U12257 ( .B1(n1300), .B2(n1331), .A(n1831), .ZN(N12962) );
  aor21d1 U12258 ( .B1(n1242), .B2(n1191), .A(n1280), .Z(n1832) );
  aoi311d1 U12259 ( .C1(n1001), .C2(n962), .C3(n1042), .A(n1832), .B(n1097), 
        .ZN(n1834) );
  aoi21d1 U12260 ( .B1(n1144), .B2(n1247), .A(n1832), .ZN(n1833) );
  nr13d1 U12261 ( .A1(n1343), .A2(n1834), .A3(n1833), .ZN(N12946) );
  nd03d0 U12262 ( .A1(n1085), .A2(n1028), .A3(n1140), .ZN(n1835) );
  oaim21d1 U12263 ( .B1(n1115), .B2(n1146), .A(n1835), .ZN(n1837) );
  aoi22d1 U12264 ( .A1(n1324), .A2(n1225), .B1(n1284), .B2(n1334), .ZN(n1836)
         );
  aoim31d1 U12265 ( .B1(n1282), .B2(n1183), .B3(n1837), .A(n1836), .ZN(N12930)
         );
  oan211d1 U12266 ( .C1(n967), .C2(n1005), .B(n1056), .A(n1098), .ZN(n1840) );
  aoi21d1 U12267 ( .B1(n1232), .B2(n1184), .A(n1309), .ZN(n1839) );
  aoi21d1 U12268 ( .B1(n1144), .B2(n1221), .A(n1832), .ZN(n1838) );
  aoi211d1 U12269 ( .C1(n1840), .C2(n1839), .A(n1351), .B(n1838), .ZN(N12914)
         );
  oai21d1 U12270 ( .B1(n1060), .B2(n1095), .A(n1146), .ZN(n1841) );
  oai321d1 U12271 ( .C1(n1843), .C2(n1276), .C3(n1187), .B1(n1236), .B2(n1290), 
        .A(n1333), .ZN(n1842) );
  aoi21d1 U12272 ( .B1(n1232), .B2(n1185), .A(n1305), .ZN(n1844) );
  oaim21d1 U12273 ( .B1(n1020), .B2(n975), .A(n1844), .ZN(n1846) );
  oaim21d1 U12274 ( .B1(n1156), .B2(n1236), .A(n1844), .ZN(n1845) );
  ora311d1 U12275 ( .C1(n1091), .C2(n1044), .C3(n1846), .A(n1845), .B(n1334), 
        .Z(N12882) );
  oai21d1 U12276 ( .B1(n1012), .B2(n1058), .A(n1146), .ZN(n1847) );
  oaim21d1 U12277 ( .B1(n1115), .B2(n1148), .A(n1847), .ZN(n1849) );
  aoi22d1 U12278 ( .A1(n1324), .A2(n1225), .B1(n1284), .B2(n1332), .ZN(n1848)
         );
  aoim31d1 U12279 ( .B1(n1282), .B2(n1184), .B3(n1849), .A(n1848), .ZN(N12866)
         );
  aoi21d1 U12280 ( .B1(n1233), .B2(n1185), .A(n1307), .ZN(n1852) );
  nr03d0 U12281 ( .A1(n1022), .A2(n1119), .A3(n1085), .ZN(n1851) );
  aoi21d1 U12282 ( .B1(n1143), .B2(n1257), .A(n1829), .ZN(n1850) );
  aoi311d1 U12283 ( .C1(n1852), .C2(n992), .C3(n1851), .A(n1360), .B(n1850), 
        .ZN(N12850) );
  oan211d1 U12284 ( .C1(n1135), .C2(n1183), .B(n1230), .A(n1275), .ZN(n1853)
         );
  oan211d1 U12285 ( .C1(n1135), .C2(n1182), .B(n1231), .A(n1276), .ZN(n1855)
         );
  nd04d0 U12286 ( .A1(n1120), .A2(n1039), .A3(n1024), .A4(n981), .ZN(n1854) );
  aoi221d1 U12287 ( .B1(n1855), .B2(n1854), .C1(n1855), .C2(n1266), .A(n1359), 
        .ZN(N12818) );
  aor31d1 U12288 ( .B1(n1069), .B2(n1016), .B3(n1093), .A(n1147), .Z(n1857) );
  aoi22d1 U12289 ( .A1(n1329), .A2(n1225), .B1(n1284), .B2(n1330), .ZN(n1856)
         );
  aoim31d1 U12290 ( .B1(n1281), .B2(n1184), .B3(n1857), .A(n1856), .ZN(N12802)
         );
  oan211d1 U12291 ( .C1(n1135), .C2(n1182), .B(n1230), .A(n1276), .ZN(n1859)
         );
  oai211d1 U12292 ( .C1(n959), .C2(n1017), .A(n1065), .B(n1095), .ZN(n1858) );
  aoi221d1 U12293 ( .B1(n1859), .B2(n1858), .C1(n1859), .C2(n1222), .A(n1359), 
        .ZN(N12786) );
  aor21d1 U12294 ( .B1(n1112), .B2(n1061), .A(n1145), .Z(n1860) );
  oai321d1 U12295 ( .C1(n1860), .C2(n1276), .C3(n1187), .B1(n1250), .B2(n1290), 
        .A(n1333), .ZN(n1861) );
  aoi321d1 U12296 ( .C1(n969), .C2(n1090), .C3(n1000), .B1(n1108), .B2(n1054), 
        .A(n2546), .ZN(n1862) );
  aoim2m11d1 U12297 ( .C1(n1883), .C2(n1227), .B(n1325), .A(n1862), .ZN(N12754) );
  oan211d1 U12298 ( .C1(n1006), .C2(n1048), .B(n1093), .A(n1141), .ZN(n1863)
         );
  aoi22d1 U12299 ( .A1(n1328), .A2(n1225), .B1(n1284), .B2(N11556), .ZN(n1864)
         );
  aoim31d1 U12300 ( .B1(n1205), .B2(n1273), .B3(n1865), .A(n1864), .ZN(N12738)
         );
  oai21d1 U12301 ( .B1(n969), .B2(n1009), .A(n1104), .ZN(n1866) );
  aoi211d1 U12302 ( .C1(n1106), .C2(n1056), .A(n2546), .B(n1868), .ZN(n1867)
         );
  aoim2m11d1 U12303 ( .C1(n1883), .C2(n1227), .B(n1342), .A(n1867), .ZN(N12722) );
  oan211d1 U12304 ( .C1(n1092), .C2(n1132), .B(n1229), .A(n1276), .ZN(n1869)
         );
  aon211d1 U12305 ( .C1(n1225), .C2(n1179), .B(n1871), .A(n1331), .ZN(n1870)
         );
  aoi311d1 U12306 ( .C1(n1001), .C2(n962), .C3(n1043), .A(n2546), .B(n1110), 
        .ZN(n1872) );
  aoim2m11d1 U12307 ( .C1(n2546), .C2(n1227), .B(n1325), .A(n1872), .ZN(N12690) );
  aoi21d1 U12308 ( .B1(n1059), .B2(n1006), .A(n1110), .ZN(n1875) );
  nr03d0 U12309 ( .A1(n1159), .A2(n1289), .A3(n1195), .ZN(n1874) );
  aoi22d1 U12310 ( .A1(n1326), .A2(n1225), .B1(n1285), .B2(n1324), .ZN(n1873)
         );
  aoi21d1 U12311 ( .B1(n1875), .B2(n1874), .A(n1873), .ZN(N12674) );
  oan211d1 U12312 ( .C1(n966), .C2(n1004), .B(n1057), .A(n1099), .ZN(n1877) );
  oan211d1 U12313 ( .C1(n1135), .C2(n1182), .B(n1230), .A(n1276), .ZN(n1876)
         );
  aoi221d1 U12314 ( .B1(n1877), .B2(n1876), .C1(n1876), .C2(n1269), .A(n1359), 
        .ZN(N12658) );
  or03d0 U12315 ( .A1(n1280), .A2(n1202), .A3(n1157), .Z(n1878) );
  oai321d1 U12316 ( .C1(n1878), .C2(n1099), .C3(n1053), .B1(n1246), .B2(n1290), 
        .A(n1333), .ZN(n1879) );
  oan211d1 U12317 ( .C1(n1135), .C2(n1182), .B(n1229), .A(n1276), .ZN(n1880)
         );
  oaim21d1 U12318 ( .B1(n1020), .B2(n975), .A(n1880), .ZN(n1881) );
  oai321d1 U12319 ( .C1(n1881), .C2(n1099), .C3(n1052), .B1(n1226), .B2(n1883), 
        .A(n1333), .ZN(n1882) );
  nr03d0 U12320 ( .A1(n1022), .A2(n1119), .A3(n1038), .ZN(n1886) );
  nr03d0 U12321 ( .A1(n1152), .A2(n1288), .A3(n1189), .ZN(n1885) );
  aoi22d1 U12322 ( .A1(n1327), .A2(n1225), .B1(n1284), .B2(n1341), .ZN(n1884)
         );
  aoi21d1 U12323 ( .B1(n1886), .B2(n1885), .A(n1884), .ZN(N12610) );
  or03d0 U12324 ( .A1(n1093), .A2(n1051), .A3(n1002), .Z(n1887) );
  oai321d1 U12325 ( .C1(n1887), .C2(n968), .C3(n1883), .B1(n1251), .B2(n2546), 
        .A(n1333), .ZN(n1888) );
  oai21d1 U12326 ( .B1(n1234), .B2(n1275), .A(n1329), .ZN(n1889) );
  nr02d0 U12327 ( .A1(n1254), .A2(n1305), .ZN(n1892) );
  nd04d0 U12328 ( .A1(n1120), .A2(n1075), .A3(n1025), .A4(n981), .ZN(n1891) );
  aoi21d1 U12329 ( .B1(n1190), .B2(n1135), .A(n1912), .ZN(n1890) );
  aoi211d1 U12330 ( .C1(n1892), .C2(n1891), .A(n1351), .B(n1890), .ZN(N12562)
         );
  an04d0 U12331 ( .A1(n1159), .A2(n1115), .A3(n1080), .A4(n1019), .Z(n1895) );
  an02d0 U12332 ( .A1(n1339), .A2(n1296), .Z(n1893) );
  oan211d1 U12333 ( .C1(n1187), .C2(n1226), .B(n1326), .A(n1893), .ZN(n1894)
         );
  aoim31d1 U12334 ( .B1(n1243), .B2(n1288), .B3(n1895), .A(n1894), .ZN(N12546)
         );
  nr02d0 U12335 ( .A1(n1254), .A2(n1306), .ZN(n1898) );
  oai211d1 U12336 ( .C1(n959), .C2(n1028), .A(n1065), .B(n1095), .ZN(n1897) );
  aoi21d1 U12337 ( .B1(n1190), .B2(n1132), .A(n2556), .ZN(n1896) );
  aoi211d1 U12338 ( .C1(n1898), .C2(n1897), .A(n1354), .B(n1896), .ZN(N12530)
         );
  an03d0 U12339 ( .A1(n1098), .A2(n1079), .A3(n1157), .Z(n1900) );
  oai21d1 U12340 ( .B1(n1279), .B2(n1231), .A(n1329), .ZN(n1899) );
  oaim31d1 U12341 ( .B1(n1334), .B2(n1193), .B3(n1900), .A(n1899), .ZN(N12514)
         );
  or02d0 U12342 ( .A1(n1234), .A2(n1302), .Z(n1901) );
  aoi21d1 U12343 ( .B1(n1190), .B2(n1161), .A(n1901), .ZN(n1903) );
  aoi321d1 U12344 ( .C1(n970), .C2(n1090), .C3(n1027), .B1(n1108), .B2(n1055), 
        .A(n1901), .ZN(n1902) );
  nr13d1 U12345 ( .A1(n1343), .A2(n1903), .A3(n1902), .ZN(N12498) );
  ora211d1 U12346 ( .C1(n1002), .C2(n1060), .A(n1116), .B(n1155), .Z(n1906) );
  an02d0 U12347 ( .A1(n1339), .A2(n1296), .Z(n1904) );
  oan211d1 U12348 ( .C1(n1187), .C2(n1248), .B(n1326), .A(n1904), .ZN(n1905)
         );
  aoim31d1 U12349 ( .B1(n1235), .B2(n1287), .B3(n1906), .A(n1905), .ZN(N12482)
         );
  oai21d1 U12350 ( .B1(n970), .B2(n1009), .A(n1105), .ZN(n1910) );
  nd02d0 U12351 ( .A1(n1095), .A2(n1083), .ZN(n1909) );
  nr02d0 U12352 ( .A1(n1255), .A2(n1305), .ZN(n1908) );
  aoi21d1 U12353 ( .B1(n1190), .B2(n1150), .A(n2578), .ZN(n1907) );
  aoi311d1 U12354 ( .C1(n1910), .C2(n1909), .C3(n1908), .A(n1359), .B(n1907), 
        .ZN(N12466) );
  aor311d1 U12355 ( .C1(n1154), .C2(n1110), .C3(n1186), .A(n1293), .B(n1253), 
        .Z(n1911) );
  an02d0 U12356 ( .A1(n1339), .A2(n1911), .Z(N12450) );
  or02d0 U12357 ( .A1(n1244), .A2(n1302), .Z(n1912) );
  aoi21d1 U12358 ( .B1(n1190), .B2(n1149), .A(n1912), .ZN(n1914) );
  aoi311d1 U12359 ( .C1(n1026), .C2(n963), .C3(n1042), .A(n1912), .B(n1109), 
        .ZN(n1913) );
  nr13d1 U12360 ( .A1(n1343), .A2(n1914), .A3(n1913), .ZN(N12434) );
  oai21d1 U12361 ( .B1(n1191), .B2(n1231), .A(n1329), .ZN(n1917) );
  nd12d0 U12362 ( .A1(n1255), .A2(n1319), .ZN(n1915) );
  aoi321d1 U12363 ( .C1(n1060), .C2(n1002), .C3(n1134), .B1(n1109), .B2(n1136), 
        .A(n1915), .ZN(n1916) );
  oan211d1 U12364 ( .C1(n1358), .C2(n1319), .B(n1917), .A(n1916), .ZN(N12418)
         );
  oan211d1 U12365 ( .C1(n966), .C2(n1004), .B(n1057), .A(n1099), .ZN(n1920) );
  nr02d0 U12366 ( .A1(n1254), .A2(n1306), .ZN(n1919) );
  aoi21d1 U12367 ( .B1(n1190), .B2(n1155), .A(n2570), .ZN(n1918) );
  aoi211d1 U12368 ( .C1(n1920), .C2(n1919), .A(n1356), .B(n1918), .ZN(N12402)
         );
  ora211d1 U12369 ( .C1(n1046), .C2(n1102), .A(n1157), .B(n1200), .Z(n1921) );
  ora31d1 U12370 ( .B1(n1277), .B2(n1238), .B3(n1921), .A(n1338), .Z(N12386)
         );
  nr02d0 U12371 ( .A1(n1255), .A2(n1306), .ZN(n1922) );
  oaim21d1 U12372 ( .B1(n1020), .B2(n983), .A(n1922), .ZN(n1924) );
  oaim21d1 U12373 ( .B1(n1201), .B2(n1148), .A(n1922), .ZN(n1923) );
  ora311d1 U12374 ( .C1(n1107), .C2(n1044), .C3(n1924), .A(n1923), .B(n1334), 
        .Z(N12370) );
  or02d0 U12375 ( .A1(n1027), .A2(n1076), .Z(n1925) );
  aor22d1 U12376 ( .A1(n1152), .A2(n1925), .B1(n1111), .B2(n1135), .Z(n1928)
         );
  an02d0 U12377 ( .A1(n1338), .A2(n1296), .Z(n1926) );
  oan211d1 U12378 ( .C1(n1187), .C2(n1255), .B(n1326), .A(n1926), .ZN(n1927)
         );
  aoim31d1 U12379 ( .B1(n1246), .B2(n1306), .B3(n1928), .A(n1927), .ZN(N12354)
         );
  nr02d0 U12380 ( .A1(n1290), .A2(n1250), .ZN(n1931) );
  nr03d0 U12381 ( .A1(n1022), .A2(n1119), .A3(n1084), .ZN(n1930) );
  aoi21d1 U12382 ( .B1(n1190), .B2(n1160), .A(n1970), .ZN(n1929) );
  aoi311d1 U12383 ( .C1(n1931), .C2(n992), .C3(n1930), .A(n1360), .B(n1929), 
        .ZN(N12338) );
  aoi211d1 U12384 ( .C1(n1198), .C2(n1138), .A(n1281), .B(n1236), .ZN(n1932)
         );
  nr02d0 U12385 ( .A1(n1932), .A2(n1370), .ZN(N12322) );
  aoi211d1 U12386 ( .C1(n1192), .C2(n1138), .A(n1281), .B(n1233), .ZN(n1934)
         );
  nd04d0 U12387 ( .A1(n1120), .A2(n1086), .A3(n1025), .A4(n982), .ZN(n1933) );
  aoi221d1 U12388 ( .B1(n1934), .B2(n1933), .C1(n1934), .C2(n1218), .A(n1359), 
        .ZN(N12306) );
  aor31d1 U12389 ( .B1(n1069), .B2(n1015), .B3(n1092), .A(n1147), .Z(n1937) );
  an02d0 U12390 ( .A1(n1339), .A2(n1295), .Z(n1935) );
  oan211d1 U12391 ( .C1(n1187), .C2(n1249), .B(n1326), .A(n1935), .ZN(n1936)
         );
  aoim31d1 U12392 ( .B1(n1229), .B2(n1300), .B3(n1937), .A(n1936), .ZN(N12290)
         );
  aoi211d1 U12393 ( .C1(n1192), .C2(n1138), .A(n1281), .B(n1242), .ZN(n1939)
         );
  oai211d1 U12394 ( .C1(n959), .C2(n1014), .A(n1066), .B(n1095), .ZN(n1938) );
  aoi221d1 U12395 ( .B1(n1939), .B2(n1938), .C1(n1939), .C2(n1219), .A(n1359), 
        .ZN(N12274) );
  nd03d0 U12396 ( .A1(n1083), .A2(n1208), .A3(n1087), .ZN(n1942) );
  nd02d0 U12397 ( .A1(n1205), .A2(n1159), .ZN(n1941) );
  oai21d1 U12398 ( .B1(n1279), .B2(n1231), .A(n1328), .ZN(n1940) );
  aon211d1 U12399 ( .C1(n1942), .C2(n1941), .B(n1357), .A(n1940), .ZN(N12258)
         );
  aor211d1 U12400 ( .C1(n1194), .C2(n1144), .A(n1285), .B(n1244), .Z(n1944) );
  aoi321d1 U12401 ( .C1(n970), .C2(num_images[3]), .C3(n1000), .B1(n1109), 
        .B2(n1054), .A(n1944), .ZN(n1943) );
  aoim2m11d1 U12402 ( .C1(n1944), .C2(n1186), .B(n1325), .A(n1943), .ZN(N12242) );
  an02d0 U12403 ( .A1(n1338), .A2(n1296), .Z(n1945) );
  oan211d1 U12404 ( .C1(n1186), .C2(n1226), .B(n1326), .A(n1945), .ZN(n1946)
         );
  aoim31d1 U12405 ( .B1(n1235), .B2(n1285), .B3(n1865), .A(n1946), .ZN(N12226)
         );
  aor211d1 U12406 ( .C1(n1195), .C2(n1148), .A(n1276), .B(n1224), .Z(n1949) );
  oai21d1 U12407 ( .B1(n970), .B2(n1008), .A(n1105), .ZN(n1947) );
  aoi211d1 U12408 ( .C1(n1106), .C2(n1057), .A(n1949), .B(n1950), .ZN(n1948)
         );
  aoim2m11d1 U12409 ( .C1(n1949), .C2(n1186), .B(n1337), .A(n1948), .ZN(N12210) );
  oai21d1 U12410 ( .B1(n1101), .B2(n1140), .A(n1202), .ZN(n1951) );
  ora31d1 U12411 ( .B1(n1272), .B2(n1230), .B3(n1952), .A(n1337), .Z(N12194)
         );
  aor211d1 U12412 ( .C1(n1194), .C2(n1159), .A(n1284), .B(n1224), .Z(n1954) );
  aoi311d1 U12413 ( .C1(n1001), .C2(n962), .C3(n1042), .A(n1954), .B(n1107), 
        .ZN(n1953) );
  aoim2m11d1 U12414 ( .C1(n1954), .C2(n1186), .B(n1324), .A(n1953), .ZN(N12178) );
  oai21d1 U12415 ( .B1(n1191), .B2(n1231), .A(n1329), .ZN(n1957) );
  or03d0 U12416 ( .A1(n1274), .A2(n1248), .A3(n1157), .Z(n1955) );
  aoi211d1 U12417 ( .C1(n1063), .C2(n1008), .A(n1955), .B(n1103), .ZN(n1956)
         );
  oan211d1 U12418 ( .C1(n1358), .C2(n1319), .B(n1957), .A(n1956), .ZN(N12162)
         );
  oan211d1 U12419 ( .C1(n966), .C2(n1005), .B(n1057), .A(n1099), .ZN(n1959) );
  aoi211d1 U12420 ( .C1(n1192), .C2(n1137), .A(n1280), .B(n1234), .ZN(n1958)
         );
  aoi221d1 U12421 ( .B1(n1959), .B2(n1958), .C1(n1958), .C2(n1176), .A(n1359), 
        .ZN(N12146) );
  oai21d1 U12422 ( .B1(n1060), .B2(n1094), .A(num_images[5]), .ZN(n1960) );
  oaim21d1 U12423 ( .B1(n1156), .B2(n1193), .A(n1960), .ZN(n1961) );
  ora31d1 U12424 ( .B1(n1286), .B2(n1231), .B3(n1961), .A(n1338), .Z(N12130)
         );
  aoi211d1 U12425 ( .C1(n1192), .C2(n1138), .A(n1280), .B(n1247), .ZN(n1962)
         );
  oaim21d1 U12426 ( .B1(n1019), .B2(N6867), .A(n1962), .ZN(n1963) );
  oai321d1 U12427 ( .C1(n1963), .C2(n1099), .C3(n1053), .B1(n1185), .B2(n13), 
        .A(n1333), .ZN(n1964) );
  oai21d1 U12428 ( .B1(n1191), .B2(n1231), .A(n1329), .ZN(n1967) );
  or03d0 U12429 ( .A1(n1278), .A2(n1226), .A3(n1157), .Z(n1965) );
  nr04d0 U12430 ( .A1(n1965), .A2(n1022), .A3(n1106), .A4(n1071), .ZN(n1966)
         );
  oan211d1 U12431 ( .C1(n1358), .C2(n1319), .B(n1967), .A(n1966), .ZN(N12098)
         );
  or02d0 U12432 ( .A1(n1276), .A2(n1248), .Z(n1970) );
  or03d0 U12433 ( .A1(n1141), .A2(n1117), .A3(n1041), .Z(n1968) );
  nr04d0 U12434 ( .A1(n1968), .A2(n1970), .A3(n1026), .A4(n979), .ZN(n1969) );
  aoim2m11d1 U12435 ( .C1(n1193), .C2(n1970), .B(n1325), .A(n1969), .ZN(N12082) );
  oai21d1 U12436 ( .B1(n1191), .B2(n1231), .A(n1329), .ZN(n1971) );
  oaim21d1 U12437 ( .B1(n1300), .B2(n1327), .A(n1971), .ZN(N12066) );
  nr03d0 U12438 ( .A1(n1307), .A2(n1248), .A3(n1197), .ZN(n1973) );
  nd04d0 U12439 ( .A1(n1120), .A2(n1072), .A3(n1024), .A4(n981), .ZN(n1972) );
  aoi22d1 U12440 ( .A1(n1973), .A2(n1972), .B1(n1171), .B2(n1973), .ZN(n1974)
         );
  an02d0 U12441 ( .A1(n1974), .A2(n1337), .Z(N12050) );
  nd04d0 U12442 ( .A1(n1162), .A2(n1104), .A3(n1075), .A4(n1023), .ZN(n1975)
         );
  nd12d0 U12443 ( .A1(num_images[5]), .A2(n1975), .ZN(n1976) );
  ora31d1 U12444 ( .B1(n1279), .B2(n1223), .B3(n1976), .A(n1338), .Z(N12034)
         );
  nr03d0 U12445 ( .A1(n1307), .A2(n1225), .A3(n1196), .ZN(n1978) );
  oai211d1 U12446 ( .C1(n959), .C2(n999), .A(n1065), .B(n1095), .ZN(n1977) );
  aoi22d1 U12447 ( .A1(n1978), .A2(n1977), .B1(n1173), .B2(n1978), .ZN(n1979)
         );
  an02d0 U12448 ( .A1(n1979), .A2(n1337), .Z(N12018) );
  aor31d1 U12449 ( .B1(n1112), .B2(n1064), .B3(n1135), .A(n1193), .Z(n1980) );
  ora31d1 U12450 ( .B1(n1298), .B2(n1223), .B3(n1980), .A(n1338), .Z(N12002)
         );
  or03d0 U12451 ( .A1(n1286), .A2(n1248), .A3(n1200), .Z(n1982) );
  aoi321d1 U12452 ( .C1(n971), .C2(n1087), .C3(n1000), .B1(n1107), .B2(n1055), 
        .A(n1982), .ZN(n1981) );
  aoim2m11d1 U12453 ( .C1(n1145), .C2(n1982), .B(n1325), .A(n1981), .ZN(N11986) );
  oai211d1 U12454 ( .C1(n998), .C2(n1043), .A(n1111), .B(n1140), .ZN(n1983) );
  nd12d0 U12455 ( .A1(num_images[5]), .A2(n1983), .ZN(n1984) );
  ora31d1 U12456 ( .B1(n1291), .B2(n1223), .B3(n1984), .A(n1338), .Z(N11970)
         );
  or03d0 U12457 ( .A1(n1281), .A2(n1254), .A3(n1198), .Z(n1987) );
  oai21d1 U12458 ( .B1(n971), .B2(n1008), .A(n1105), .ZN(n1985) );
  aoi211d1 U12459 ( .C1(n1106), .C2(n1057), .A(n1987), .B(n1988), .ZN(n1986)
         );
  aoim2m11d1 U12460 ( .C1(n1146), .C2(n1987), .B(n1325), .A(n1986), .ZN(N11954) );
  aor21d1 U12461 ( .B1(n1137), .B2(n1101), .A(n1180), .Z(n1989) );
  ora31d1 U12462 ( .B1(n1294), .B2(n1223), .B3(n1989), .A(n1338), .Z(N11938)
         );
  or03d0 U12463 ( .A1(n1275), .A2(n1248), .A3(n1199), .Z(n1991) );
  aoi311d1 U12464 ( .C1(n1001), .C2(n962), .C3(n1043), .A(n1991), .B(n1108), 
        .ZN(n1990) );
  aoim2m11d1 U12465 ( .C1(n1145), .C2(n1991), .B(n1325), .A(n1990), .ZN(N11922) );
  nd02d0 U12466 ( .A1(n1118), .A2(n1159), .ZN(n1994) );
  nd03d0 U12467 ( .A1(n1081), .A2(n1028), .A3(n1154), .ZN(n1993) );
  nr03d0 U12468 ( .A1(n1203), .A2(n1290), .A3(n1225), .ZN(n1992) );
  aoi31d1 U12469 ( .B1(n1994), .B2(n1993), .B3(n1992), .A(n1366), .ZN(N11906)
         );
  oan211d1 U12470 ( .C1(n965), .C2(n1004), .B(n1056), .A(n1099), .ZN(n1996) );
  nr03d0 U12471 ( .A1(n1307), .A2(n1230), .A3(n1202), .ZN(n1995) );
  aoi22d1 U12472 ( .A1(n1996), .A2(n1995), .B1(n1174), .B2(n1995), .ZN(n1997)
         );
  an02d0 U12473 ( .A1(n1997), .A2(n1337), .Z(N11890) );
  oan211d1 U12474 ( .C1(n1051), .C2(n1094), .B(n1138), .A(n1189), .ZN(n1998)
         );
  ora31d1 U12475 ( .B1(n1297), .B2(n1223), .B3(n1999), .A(n1337), .Z(N11874)
         );
  nr03d0 U12476 ( .A1(n1307), .A2(n1250), .A3(n1193), .ZN(n2000) );
  oaim21d1 U12477 ( .B1(n1019), .B2(n957), .A(n2000), .ZN(n2001) );
  oai321d1 U12478 ( .C1(n2001), .C2(n1099), .C3(n1052), .B1(n1135), .B2(n8), 
        .A(n1334), .ZN(n2002) );
  nd02d0 U12479 ( .A1(n1107), .A2(n1159), .ZN(n2005) );
  oai21d1 U12480 ( .B1(n1013), .B2(n1058), .A(n1146), .ZN(n2004) );
  nr03d0 U12481 ( .A1(n1202), .A2(n1305), .A3(n1245), .ZN(n2003) );
  aoi31d1 U12482 ( .B1(n2005), .B2(n2004), .B3(n2003), .A(n1366), .ZN(N11842)
         );
  nr02d0 U12483 ( .A1(n1303), .A2(n1250), .ZN(n2007) );
  nr02d0 U12484 ( .A1(n1026), .A2(n978), .ZN(n2008) );
  nr03d0 U12485 ( .A1(n1070), .A2(n1206), .A3(n1119), .ZN(n2006) );
  nd03d0 U12486 ( .A1(n2008), .A2(n2007), .A3(n2006), .ZN(n2009) );
  ora311d1 U12487 ( .C1(n1183), .C2(n1142), .C3(n1970), .A(n2009), .B(n1334), 
        .Z(N11826) );
  nr04d0 U12488 ( .A1(n1304), .A2(n1252), .A3(n1175), .A4(n1161), .ZN(n2010)
         );
  nr02d0 U12489 ( .A1(n2010), .A2(n1369), .ZN(N11810) );
  nd04d0 U12490 ( .A1(n1110), .A2(n1072), .A3(n1025), .A4(n982), .ZN(n2012) );
  nr03d0 U12491 ( .A1(n1203), .A2(n1277), .A3(n1230), .ZN(n2011) );
  aoi31d1 U12492 ( .B1(n2012), .B2(n1171), .B3(n2011), .A(n1366), .ZN(N11794)
         );
  aoi31d1 U12493 ( .B1(n1068), .B2(n1005), .B3(n1107), .A(n1149), .ZN(n2014)
         );
  nr03d0 U12494 ( .A1(n1203), .A2(n1306), .A3(n1226), .ZN(n2013) );
  aoi21d1 U12495 ( .B1(n2014), .B2(n2013), .A(n1356), .ZN(N11778) );
  oai211d1 U12496 ( .C1(n998), .C2(n961), .A(n1065), .B(n1095), .ZN(n2016) );
  nr03d0 U12497 ( .A1(n1202), .A2(n1301), .A3(n1233), .ZN(n2015) );
  aoi31d1 U12498 ( .B1(n2016), .B2(n1171), .B3(n2015), .A(n1371), .ZN(N11762)
         );
  aoi21d1 U12499 ( .B1(n1101), .B2(n1049), .A(n1155), .ZN(n2018) );
  nr03d0 U12500 ( .A1(n1203), .A2(n1304), .A3(n1232), .ZN(n2017) );
  aoi21d1 U12501 ( .B1(n2018), .B2(n2017), .A(n1368), .ZN(N11746) );
  aoi321d1 U12502 ( .C1(n971), .C2(n1091), .C3(n1026), .B1(n1107), .B2(n1055), 
        .A(n1155), .ZN(n2020) );
  nr03d0 U12503 ( .A1(n1203), .A2(num_images[7]), .A3(n1223), .ZN(n2019) );
  aoi21d1 U12504 ( .B1(n2020), .B2(n2019), .A(n1367), .ZN(N11730) );
  oan211d1 U12505 ( .C1(n1007), .C2(n1048), .B(n1093), .A(n1140), .ZN(n2022)
         );
  nr03d0 U12506 ( .A1(n1203), .A2(n1272), .A3(n1255), .ZN(n2021) );
  aoi21d1 U12507 ( .B1(n2022), .B2(n2021), .A(n1370), .ZN(N11714) );
  aoi21d1 U12508 ( .B1(n1101), .B2(n1049), .A(n1150), .ZN(n2025) );
  oai21d1 U12509 ( .B1(n1013), .B2(n968), .A(n1104), .ZN(n2024) );
  nr03d0 U12510 ( .A1(n1203), .A2(n1307), .A3(n1224), .ZN(n2023) );
  aoi31d1 U12511 ( .B1(n2025), .B2(n2024), .B3(n2023), .A(n1369), .ZN(N11698)
         );
  or03d0 U12512 ( .A1(n1293), .A2(n1248), .A3(n1196), .Z(n2026) );
  ora31d1 U12513 ( .B1(n1157), .B2(n1089), .B3(n2026), .A(n1337), .Z(N11682)
         );
  aoi311d1 U12514 ( .C1(num_images[1]), .C2(n962), .C3(n1042), .A(n1137), .B(
        n1115), .ZN(n2028) );
  nr03d0 U12515 ( .A1(n1203), .A2(n1302), .A3(n1230), .ZN(n2027) );
  aoi21d1 U12516 ( .B1(n2028), .B2(n2027), .A(n1372), .ZN(N11666) );
  aoi211d1 U12517 ( .C1(n1062), .C2(n1008), .A(n1146), .B(n1089), .ZN(n2030)
         );
  nr03d0 U12518 ( .A1(n1203), .A2(n1273), .A3(n1228), .ZN(n2029) );
  aoi21d1 U12519 ( .B1(n2030), .B2(n2029), .A(n1366), .ZN(N11650) );
  nr02d0 U12520 ( .A1(n1162), .A2(n1118), .ZN(n2033) );
  oai21d1 U12521 ( .B1(n1013), .B2(n968), .A(n1062), .ZN(n2032) );
  nr03d0 U12522 ( .A1(n1203), .A2(n1287), .A3(n1248), .ZN(n2031) );
  aoi31d1 U12523 ( .B1(n2033), .B2(n2032), .B3(n2031), .A(n1371), .ZN(N11634)
         );
  nr03d0 U12524 ( .A1(n1070), .A2(n1142), .A3(n1115), .ZN(n2035) );
  nr03d0 U12525 ( .A1(n1203), .A2(n1282), .A3(n1225), .ZN(n2034) );
  aoi21d1 U12526 ( .B1(n2035), .B2(n2034), .A(n1367), .ZN(N11618) );
  aoi211d1 U12527 ( .C1(n1014), .C2(n967), .A(n1102), .B(n1045), .ZN(n2037) );
  nr04d0 U12528 ( .A1(n1303), .A2(n1252), .A3(n1175), .A4(n1161), .ZN(n2036)
         );
  aoi21d1 U12529 ( .B1(n2037), .B2(n2036), .A(n1365), .ZN(N11602) );
  nr03d0 U12530 ( .A1(n1022), .A2(n1119), .A3(n1039), .ZN(n2039) );
  nr04d0 U12531 ( .A1(n1303), .A2(n1252), .A3(n1175), .A4(n1161), .ZN(n2038)
         );
  aoi21d1 U12532 ( .B1(n2039), .B2(n2038), .A(n1365), .ZN(N11586) );
  nr04d0 U12533 ( .A1(n1092), .A2(n1070), .A3(n1027), .A4(n979), .ZN(n2041) );
  nr04d0 U12534 ( .A1(n1303), .A2(n1252), .A3(n1175), .A4(n1148), .ZN(n2040)
         );
  aoi21d1 U12535 ( .B1(n2041), .B2(n2040), .A(n1365), .ZN(N11571) );
  nd04d0 U12536 ( .A1(n1094), .A2(n1072), .A3(n1026), .A4(n981), .ZN(n2043) );
  nd04d0 U12537 ( .A1(n1305), .A2(n1256), .A3(n1207), .A4(n1154), .ZN(n2042)
         );
  oai21d1 U12538 ( .B1(n2043), .B2(n2042), .A(n1361), .ZN(N11541) );
  nd04d0 U12539 ( .A1(n1162), .A2(n1106), .A3(n1076), .A4(n1023), .ZN(n2045)
         );
  aoi31d1 U12540 ( .B1(n1239), .B2(n1194), .B3(n1286), .A(n1342), .ZN(n2044)
         );
  aoi21d1 U12541 ( .B1(n2045), .B2(n1357), .A(n2044), .ZN(N11526) );
  nd03d0 U12542 ( .A1(n1239), .A2(n1209), .A3(n1276), .ZN(n2048) );
  oai21d1 U12543 ( .B1(n1013), .B2(n968), .A(n1062), .ZN(n2047) );
  nd02d0 U12544 ( .A1(n1161), .A2(n1100), .ZN(n2046) );
  oai31d1 U12545 ( .B1(n2048), .B2(n2047), .B3(n2046), .A(n1369), .ZN(N11511)
         );
  nd04d0 U12546 ( .A1(n1200), .A2(n1141), .A3(n1106), .A4(n1071), .ZN(n2050)
         );
  aoi21d1 U12547 ( .B1(n1278), .B2(num_images[6]), .A(n1344), .ZN(n2049) );
  aoi21d1 U12548 ( .B1(n2050), .B2(n1358), .A(n2049), .ZN(N11496) );
  nd03d0 U12549 ( .A1(n1001), .A2(n983), .A3(n1097), .ZN(n2051) );
  oaim21d1 U12550 ( .B1(n1076), .B2(n1098), .A(n2051), .ZN(n2052) );
  an03d0 U12551 ( .A1(n1161), .A2(n2052), .A3(n1201), .Z(n2053) );
  aor31d1 U12552 ( .B1(n1294), .B2(n1237), .B3(n2053), .A(n1330), .Z(N11481)
         );
  oai211d1 U12553 ( .C1(n998), .C2(n1043), .A(n1110), .B(n1139), .ZN(n2055) );
  aoi31d1 U12554 ( .B1(n1239), .B2(n1194), .B3(n1286), .A(n1332), .ZN(n2054)
         );
  aoi21d1 U12555 ( .B1(n2055), .B2(n1358), .A(n2054), .ZN(N11466) );
  ora311d1 U12556 ( .C1(n1046), .C2(num_images[1]), .C3(n963), .A(n1114), .B(
        n1154), .Z(n2056) );
  nd04d0 U12557 ( .A1(n1255), .A2(n1208), .A3(n1296), .A4(n2056), .ZN(n2057)
         );
  nd12d0 U12558 ( .A1(n1349), .A2(n2057), .ZN(N11451) );
  nd04d0 U12559 ( .A1(n1255), .A2(n1208), .A3(n1135), .A4(n1114), .ZN(n2058)
         );
  aoim22d1 U12560 ( .A1(n2058), .A2(n1357), .B1(n1293), .B2(n1332), .Z(N11436)
         );
  aor31d1 U12561 ( .B1(n1018), .B2(n977), .B3(n1052), .A(n1106), .Z(n2059) );
  an03d0 U12562 ( .A1(n1161), .A2(n2059), .A3(n1185), .Z(n2060) );
  aor31d1 U12563 ( .B1(n1294), .B2(n1237), .B3(n2060), .A(n1330), .Z(N11421)
         );
  nd03d0 U12564 ( .A1(n1254), .A2(n1209), .A3(n1300), .ZN(n2062) );
  aoi321d1 U12565 ( .C1(n1059), .C2(n1003), .C3(n1134), .B1(n1108), .B2(n1136), 
        .A(n1336), .ZN(n2061) );
  aoi21d1 U12566 ( .B1(n2062), .B2(n1358), .A(n2061), .ZN(N11406) );
  oai321d1 U12567 ( .C1(n965), .C2(n1098), .C3(n1008), .B1(n1090), .B2(n1063), 
        .A(n1140), .ZN(n2064) );
  nd03d0 U12568 ( .A1(n1227), .A2(n1209), .A3(n1270), .ZN(n2063) );
  oai21d1 U12569 ( .B1(n2064), .B2(n2063), .A(n1361), .ZN(N11391) );
  oai211d1 U12570 ( .C1(n1042), .C2(n1090), .A(n1153), .B(n1189), .ZN(n2066)
         );
  aoi21d1 U12571 ( .B1(n1278), .B2(num_images[6]), .A(n1338), .ZN(n2065) );
  aoi21d1 U12572 ( .B1(n2066), .B2(n1358), .A(n2065), .ZN(N11376) );
  aor211d1 U12573 ( .C1(n1016), .C2(n964), .A(n1089), .B(n1046), .Z(n2067) );
  an03d0 U12574 ( .A1(n1161), .A2(n1190), .A3(n2067), .Z(n2068) );
  oan211d1 U12575 ( .C1(n1006), .C2(n1048), .B(n1138), .A(n1328), .ZN(n2070)
         );
  aoi31d1 U12576 ( .B1(n1239), .B2(n1194), .B3(n1286), .A(n1332), .ZN(n2069)
         );
  oan211d1 U12577 ( .C1(n1133), .C2(n1128), .B(n2070), .A(n2069), .ZN(N11346)
         );
  or04d0 U12578 ( .A1(n1101), .A2(n1057), .A3(n1003), .A4(n983), .Z(n2071) );
  an03d0 U12579 ( .A1(n1161), .A2(n1179), .A3(n2071), .Z(n2072) );
  aor31d1 U12580 ( .B1(n1294), .B2(n1237), .B3(n2072), .A(n1330), .Z(N11331)
         );
  nd04d0 U12581 ( .A1(n1291), .A2(n1256), .A3(n1207), .A4(n1136), .ZN(n2073)
         );
  nd12d0 U12582 ( .A1(n1349), .A2(n2073), .ZN(N11316) );
  nd04d0 U12583 ( .A1(n1089), .A2(n1072), .A3(n1025), .A4(n981), .ZN(n2074) );
  nd12d0 U12584 ( .A1(n1163), .A2(n2074), .ZN(n2075) );
  nd04d0 U12585 ( .A1(n1199), .A2(n1278), .A3(n1254), .A4(n2075), .ZN(n2076)
         );
  nd12d0 U12586 ( .A1(n1347), .A2(n2076), .ZN(N11301) );
  nd03d0 U12587 ( .A1(n1242), .A2(n1209), .A3(n1270), .ZN(n2078) );
  aoi311d1 U12588 ( .C1(n1045), .C2(n1028), .C3(n1116), .A(n1325), .B(n1161), 
        .ZN(n2077) );
  aoi21d1 U12589 ( .B1(n2078), .B2(n1358), .A(n2077), .ZN(N11286) );
  oai211d1 U12590 ( .C1(n959), .C2(n1021), .A(n1066), .B(n1095), .ZN(n2079) );
  nd12d0 U12591 ( .A1(n1162), .A2(n2079), .ZN(n2080) );
  nd04d0 U12592 ( .A1(num_images[5]), .A2(n1275), .A3(n1254), .A4(n2080), .ZN(
        n2081) );
  nd12d0 U12593 ( .A1(n1346), .A2(n2081), .ZN(N11271) );
  nd03d0 U12594 ( .A1(n1071), .A2(n1209), .A3(n1098), .ZN(n2082) );
  oaim21d1 U12595 ( .B1(n1201), .B2(n1141), .A(n2082), .ZN(n2083) );
  aor31d1 U12596 ( .B1(n1241), .B2(n2083), .B3(n1274), .A(n1331), .Z(N11256)
         );
  aoi321d1 U12597 ( .C1(n972), .C2(n1087), .C3(num_images[1]), .B1(n1109), 
        .B2(n1053), .A(n1155), .ZN(n2084) );
  nr02d0 U12598 ( .A1(n2084), .A2(n1222), .ZN(n2085) );
  aor31d1 U12599 ( .B1(n1198), .B2(n1291), .B3(n2085), .A(n1331), .Z(N11241)
         );
  oai21d1 U12600 ( .B1(n1013), .B2(n1058), .A(n1103), .ZN(n2086) );
  aoi31d1 U12601 ( .B1(n1239), .B2(n1200), .B3(n1286), .A(n1332), .ZN(n2087)
         );
  aoim31d1 U12602 ( .B1(n1147), .B2(n1324), .B3(n2088), .A(n2087), .ZN(N11226)
         );
  aoi21d1 U12603 ( .B1(n1100), .B2(n1050), .A(n1149), .ZN(n2090) );
  oai21d1 U12604 ( .B1(n973), .B2(n1009), .A(n1103), .ZN(n2089) );
  aoi21d1 U12605 ( .B1(n2090), .B2(n2089), .A(n1258), .ZN(n2091) );
  aor31d1 U12606 ( .B1(n1198), .B2(n1291), .B3(n2091), .A(n1331), .Z(N11211)
         );
  oai211d1 U12607 ( .C1(n1095), .C2(n1152), .A(n1189), .B(n1231), .ZN(n2092)
         );
  aoim22d1 U12608 ( .A1(n2092), .A2(n1357), .B1(n1294), .B2(n1332), .Z(N11196)
         );
  aor311d1 U12609 ( .C1(n1017), .C2(n976), .C3(n1051), .A(n1162), .B(n1104), 
        .Z(n2093) );
  nd04d0 U12610 ( .A1(num_images[5]), .A2(n1281), .A3(n1254), .A4(n2093), .ZN(
        n2094) );
  nd12d0 U12611 ( .A1(n1349), .A2(n2094), .ZN(N11181) );
  aor21d1 U12612 ( .B1(n1069), .B2(n1013), .A(n1102), .Z(n2096) );
  aoi31d1 U12613 ( .B1(n1240), .B2(n1194), .B3(n1286), .A(n1332), .ZN(n2095)
         );
  aoim31d1 U12614 ( .B1(n1147), .B2(n1324), .B3(n2096), .A(n2095), .ZN(N11166)
         );
  oai21d1 U12615 ( .B1(n972), .B2(n1008), .A(n1062), .ZN(n2097) );
  ora31d1 U12616 ( .B1(n1145), .B2(n1089), .B3(n2099), .A(n1243), .Z(n2098) );
  aor31d1 U12617 ( .B1(n1198), .B2(n1291), .B3(n2098), .A(n1331), .Z(N11151)
         );
  oan211d1 U12618 ( .C1(n1052), .C2(n1087), .B(n1188), .A(n1328), .ZN(n2101)
         );
  aoi21d1 U12619 ( .B1(n1278), .B2(n1221), .A(n1332), .ZN(n2100) );
  oan211d1 U12620 ( .C1(n1176), .C2(n1172), .B(n2101), .A(n2100), .ZN(N11136)
         );
  aor21d1 U12621 ( .B1(n1018), .B2(n972), .A(n1061), .Z(n2102) );
  ora31d1 U12622 ( .B1(n1139), .B2(n1089), .B3(n2102), .A(n1243), .Z(n2103) );
  aor31d1 U12623 ( .B1(n1198), .B2(n1291), .B3(n2103), .A(n1331), .Z(N11121)
         );
  or03d0 U12624 ( .A1(n1348), .A2(n1158), .A3(n1116), .Z(n2105) );
  aoi31d1 U12625 ( .B1(n1239), .B2(n1194), .B3(n1286), .A(n1332), .ZN(n2104)
         );
  aoim31d1 U12626 ( .B1(n1061), .B2(n1005), .B3(n2105), .A(n2104), .ZN(N11106)
         );
  or03d0 U12627 ( .A1(n1138), .A2(n1117), .A3(n1078), .Z(n2106) );
  ora31d1 U12628 ( .B1(num_images[1]), .B2(n963), .B3(n2106), .A(n1243), .Z(
        n2107) );
  aor31d1 U12629 ( .B1(n1199), .B2(n1291), .B3(n2107), .A(n1330), .Z(N11091)
         );
  aor31d1 U12630 ( .B1(n1241), .B2(n1194), .B3(n1274), .A(n1330), .Z(N11076)
         );
  an02d0 U12631 ( .A1(n1298), .A2(n1242), .Z(n2108) );
  nd02d0 U12632 ( .A1(n1205), .A2(n2108), .ZN(n2111) );
  nd04d0 U12633 ( .A1(n1099), .A2(n1072), .A3(n1025), .A4(n981), .ZN(n2110) );
  aoi21d1 U12634 ( .B1(n1143), .B2(n2108), .A(n2112), .ZN(n2109) );
  aon211d1 U12635 ( .C1(n2111), .C2(n2110), .B(n2109), .A(n1361), .ZN(N11061)
         );
  nd03d0 U12636 ( .A1(n1277), .A2(n1257), .A3(n1028), .ZN(n2115) );
  nd03d0 U12637 ( .A1(n1113), .A2(n1073), .A3(n1162), .ZN(n2114) );
  aoi31d1 U12638 ( .B1(n1239), .B2(n1194), .B3(n1286), .A(n1346), .ZN(n2113)
         );
  oai21d1 U12639 ( .B1(n2115), .B2(n2114), .A(n2113), .ZN(N11046) );
  an02d0 U12640 ( .A1(n1298), .A2(n1242), .Z(n2116) );
  nd02d0 U12641 ( .A1(n1205), .A2(n2116), .ZN(n2119) );
  oai211d1 U12642 ( .C1(n959), .C2(n999), .A(n1066), .B(n1096), .ZN(n2118) );
  aoi21d1 U12643 ( .B1(n1141), .B2(n2116), .A(n2120), .ZN(n2117) );
  aon211d1 U12644 ( .C1(n2119), .C2(n2118), .B(n2117), .A(n1362), .ZN(N11031)
         );
  nd02d0 U12645 ( .A1(n1309), .A2(n1249), .ZN(n2122) );
  aoi311d1 U12646 ( .C1(n1089), .C2(n1044), .C3(n1140), .A(n1325), .B(n1185), 
        .ZN(n2121) );
  aoi21d1 U12647 ( .B1(n2122), .B2(n1357), .A(n2121), .ZN(N11016) );
  an02d0 U12648 ( .A1(n1298), .A2(n1242), .Z(n2123) );
  nd02d0 U12649 ( .A1(n1205), .A2(n2123), .ZN(n2126) );
  nd02d0 U12650 ( .A1(n1161), .A2(n2123), .ZN(n2125) );
  aoi321d1 U12651 ( .C1(n973), .C2(n1091), .C3(num_images[1]), .B1(n1109), 
        .B2(n1053), .A(n2127), .ZN(n2124) );
  aon211d1 U12652 ( .C1(n2126), .C2(n2125), .B(n2124), .A(n1362), .ZN(N11001)
         );
  ora211d1 U12653 ( .C1(n1002), .C2(n1059), .A(n1116), .B(n1155), .Z(n2129) );
  aoi21d1 U12654 ( .B1(n1278), .B2(n1257), .A(n1332), .ZN(n2128) );
  aoim31d1 U12655 ( .B1(n1179), .B2(n1332), .B3(n2129), .A(n2128), .ZN(N10986)
         );
  an02d0 U12656 ( .A1(n1298), .A2(n1242), .Z(n2131) );
  an02d0 U12657 ( .A1(n1200), .A2(n2131), .Z(n2130) );
  aoi21d1 U12658 ( .B1(n1100), .B2(n1050), .A(n2130), .ZN(n2134) );
  oai21d1 U12659 ( .B1(n973), .B2(n1008), .A(n1103), .ZN(n2133) );
  aoi21d1 U12660 ( .B1(n1142), .B2(n2131), .A(n2130), .ZN(n2132) );
  aon211d1 U12661 ( .C1(n2134), .C2(n2133), .B(n2132), .A(n1361), .ZN(N10971)
         );
  an03d0 U12662 ( .A1(n1118), .A2(n1247), .A3(n1156), .Z(n2135) );
  aon211d1 U12663 ( .C1(n1225), .C2(n1179), .B(n2135), .A(n1278), .ZN(n2136)
         );
  nd12d0 U12664 ( .A1(n1349), .A2(n2136), .ZN(N10956) );
  an02d0 U12665 ( .A1(n1298), .A2(n1242), .Z(n2139) );
  an02d0 U12666 ( .A1(n1200), .A2(n2139), .Z(n2138) );
  aor311d1 U12667 ( .C1(n1016), .C2(n975), .C3(n1051), .A(n1092), .B(n2138), 
        .Z(n2137) );
  aon211d1 U12668 ( .C1(n1151), .C2(n2139), .B(n2138), .A(n2137), .ZN(n2140)
         );
  nd12d0 U12669 ( .A1(n1349), .A2(n2140), .ZN(N10941) );
  nd03d0 U12670 ( .A1(n1084), .A2(n1028), .A3(n1157), .ZN(n2141) );
  oaim21d1 U12671 ( .B1(n1115), .B2(n1149), .A(n2141), .ZN(n2143) );
  aoi21d1 U12672 ( .B1(n1278), .B2(num_images[6]), .A(n1331), .ZN(n2142) );
  aoim31d1 U12673 ( .B1(n1329), .B2(n1183), .B3(n2143), .A(n2142), .ZN(N10926)
         );
  an02d0 U12674 ( .A1(n1297), .A2(n1242), .Z(n2145) );
  an02d0 U12675 ( .A1(n1200), .A2(n2145), .Z(n2144) );
  nr02d0 U12676 ( .A1(n1093), .A2(n2144), .ZN(n2148) );
  oai21d1 U12677 ( .B1(n973), .B2(n1009), .A(n1062), .ZN(n2147) );
  aoi21d1 U12678 ( .B1(n1142), .B2(n2145), .A(n2144), .ZN(n2146) );
  aon211d1 U12679 ( .C1(n2148), .C2(n2147), .B(n2146), .A(n1362), .ZN(N10911)
         );
  oai21d1 U12680 ( .B1(n1059), .B2(n1096), .A(n1146), .ZN(n2149) );
  aoi21d1 U12681 ( .B1(n1277), .B2(n1227), .A(n1337), .ZN(n2150) );
  aoim31d1 U12682 ( .B1(n1201), .B2(n1324), .B3(n2151), .A(n2150), .ZN(N10896)
         );
  an02d0 U12683 ( .A1(n1297), .A2(n1242), .Z(n2153) );
  an02d0 U12684 ( .A1(n1200), .A2(n2153), .Z(n2152) );
  aoi21d1 U12685 ( .B1(n1012), .B2(n964), .A(n2152), .ZN(n2156) );
  nr02d0 U12686 ( .A1(n1115), .A2(n1041), .ZN(n2155) );
  aoi21d1 U12687 ( .B1(n1141), .B2(n2153), .A(n2152), .ZN(n2154) );
  aon211d1 U12688 ( .C1(n2156), .C2(n2155), .B(n2154), .A(n1364), .ZN(N10881)
         );
  oai21d1 U12689 ( .B1(n1012), .B2(n1058), .A(n1146), .ZN(n2157) );
  oaim21d1 U12690 ( .B1(n1115), .B2(n1135), .A(n2157), .ZN(n2159) );
  aoi21d1 U12691 ( .B1(n1277), .B2(num_images[6]), .A(n1330), .ZN(n2158) );
  aoim31d1 U12692 ( .B1(n1328), .B2(n1183), .B3(n2159), .A(n2158), .ZN(N10866)
         );
  an02d0 U12693 ( .A1(n1297), .A2(n1242), .Z(n2162) );
  or04d0 U12694 ( .A1(n1021), .A2(n977), .A3(n1097), .A4(n1062), .Z(n2160) );
  aoi31d1 U12695 ( .B1(n2162), .B2(n2160), .B3(n1148), .A(n1332), .ZN(n2161)
         );
  oaim21d1 U12696 ( .B1(n1201), .B2(n2162), .A(n2161), .ZN(N10851) );
  oai211d1 U12697 ( .C1(n1150), .C2(n1186), .A(n1238), .B(n1275), .ZN(n2163)
         );
  nd12d0 U12698 ( .A1(n1349), .A2(n2163), .ZN(N10836) );
  an02d0 U12699 ( .A1(n1019), .A2(n978), .Z(n2164) );
  aor311d1 U12700 ( .C1(n1112), .C2(n1064), .C3(n2164), .A(n1186), .B(n1134), 
        .Z(n2165) );
  aor31d1 U12701 ( .B1(n1241), .B2(n2165), .B3(n1274), .A(n1330), .Z(N10821)
         );
  aor31d1 U12702 ( .B1(n1069), .B2(n1016), .B3(n1093), .A(n1147), .Z(n2167) );
  aoi21d1 U12703 ( .B1(n1278), .B2(n1227), .A(n1343), .ZN(n2166) );
  aoim31d1 U12704 ( .B1(n1329), .B2(n1183), .B3(n2167), .A(n2166), .ZN(N10806)
         );
  or02d0 U12705 ( .A1(n983), .A2(n1021), .Z(n2168) );
  aor311d1 U12706 ( .C1(n1058), .C2(n2168), .C3(n1092), .A(n1194), .B(n1134), 
        .Z(n2169) );
  aor31d1 U12707 ( .B1(n1240), .B2(n2169), .B3(n1274), .A(n1330), .Z(N10791)
         );
  aor21d1 U12708 ( .B1(n1112), .B2(n1059), .A(n1145), .Z(n2171) );
  aoi21d1 U12709 ( .B1(n1278), .B2(n1227), .A(n1345), .ZN(n2170) );
  aoim31d1 U12710 ( .B1(n1194), .B2(n1350), .B3(n2171), .A(n2170), .ZN(N10776)
         );
  nd03d0 U12711 ( .A1(n982), .A2(n1101), .A3(n1028), .ZN(n2172) );
  oaim21d1 U12712 ( .B1(n1115), .B2(n1063), .A(n2172), .ZN(n2173) );
  oai311d1 U12713 ( .C1(n2173), .C2(n1180), .C3(n1151), .A(n1244), .B(n1293), 
        .ZN(n2174) );
  nd12d0 U12714 ( .A1(n1349), .A2(n2174), .ZN(N10761) );
  aoi21d1 U12715 ( .B1(n1278), .B2(n1227), .A(n1340), .ZN(n2175) );
  aoim31d1 U12716 ( .B1(n1179), .B2(n1341), .B3(n1865), .A(n2175), .ZN(N10746)
         );
  oai21d1 U12717 ( .B1(n974), .B2(n1009), .A(n1103), .ZN(n2177) );
  nr02d0 U12718 ( .A1(n1196), .A2(n1159), .ZN(n2176) );
  oaim211d1 U12719 ( .C1(n1113), .C2(n1067), .A(n2177), .B(n2176), .ZN(n2178)
         );
  aor31d1 U12720 ( .B1(n1241), .B2(n2178), .B3(n1274), .A(n1330), .Z(N10731)
         );
  oan211d1 U12721 ( .C1(n1093), .C2(num_images[4]), .B(n1230), .A(n1328), .ZN(
        n2180) );
  nd02d0 U12722 ( .A1(n1205), .A2(n1245), .ZN(n2179) );
  aoim22d1 U12723 ( .A1(n2180), .A2(n2179), .B1(n1294), .B2(n1333), .Z(N10716)
         );
  aor31d1 U12724 ( .B1(n1018), .B2(n977), .B3(n1052), .A(n1106), .Z(n2181) );
  oai311d1 U12725 ( .C1(n2181), .C2(n1183), .C3(n1150), .A(n1244), .B(n1293), 
        .ZN(n2182) );
  nd12d0 U12726 ( .A1(n1350), .A2(n2182), .ZN(N10701) );
  aoi21d1 U12727 ( .B1(n1058), .B2(n1005), .A(n1110), .ZN(n2185) );
  nr03d0 U12728 ( .A1(n1139), .A2(n1345), .A3(n1175), .ZN(n2184) );
  nd02d0 U12729 ( .A1(n1309), .A2(n1249), .ZN(n2183) );
  aoi22d1 U12730 ( .A1(n2185), .A2(n2184), .B1(n2183), .B2(n1357), .ZN(N10686)
         );
  oan211d1 U12731 ( .C1(n966), .C2(n1004), .B(n1055), .A(n1097), .ZN(n2187) );
  nr02d0 U12732 ( .A1(n1197), .A2(n1160), .ZN(n2186) );
  nd02d0 U12733 ( .A1(n2187), .A2(n2186), .ZN(n2188) );
  aor31d1 U12734 ( .B1(n1240), .B2(n2188), .B3(n1274), .A(n1330), .Z(N10671)
         );
  or03d0 U12735 ( .A1(n1348), .A2(n1202), .A3(n1136), .Z(n2190) );
  aoi21d1 U12736 ( .B1(n1278), .B2(n1227), .A(n1347), .ZN(n2189) );
  aoim31d1 U12737 ( .B1(n1103), .B2(n1049), .B3(n2190), .A(n2189), .ZN(N10656)
         );
  aoi21d1 U12738 ( .B1(n1012), .B2(n964), .A(n1063), .ZN(n2192) );
  nr03d0 U12739 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n2191) );
  nd02d0 U12740 ( .A1(n2192), .A2(n2191), .ZN(n2193) );
  aor31d1 U12741 ( .B1(n1241), .B2(n2193), .B3(n1274), .A(n1330), .Z(N10641)
         );
  nr03d0 U12742 ( .A1(n1022), .A2(n1119), .A3(n1074), .ZN(n2196) );
  nr03d0 U12743 ( .A1(n1160), .A2(n1346), .A3(n1191), .ZN(n2195) );
  nd02d0 U12744 ( .A1(n1303), .A2(n1249), .ZN(n2194) );
  aoi22d1 U12745 ( .A1(n2196), .A2(n2195), .B1(n2194), .B2(n1357), .ZN(N10626)
         );
  nr04d0 U12746 ( .A1(n1117), .A2(n1070), .A3(n1026), .A4(n979), .ZN(n2199) );
  nd02d0 U12747 ( .A1(n1308), .A2(n1249), .ZN(n2198) );
  oai21d1 U12748 ( .B1(n1191), .B2(n1139), .A(n1496), .ZN(n2197) );
  oai211d1 U12749 ( .C1(n2199), .C2(n2198), .A(n1368), .B(n2197), .ZN(N10611)
         );
  aor21d1 U12750 ( .B1(n1295), .B2(n1234), .A(n1328), .Z(N10596) );
  nd02d0 U12751 ( .A1(n1309), .A2(n1249), .ZN(n2202) );
  nd04d0 U12752 ( .A1(n1111), .A2(n1072), .A3(n1025), .A4(n980), .ZN(n2201) );
  aoi31d1 U12753 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n2108), .ZN(n2200)
         );
  aon211d1 U12754 ( .C1(n2202), .C2(n2201), .B(n2200), .A(n1362), .ZN(N10581)
         );
  an04d0 U12755 ( .A1(n1158), .A2(n1114), .A3(n1037), .A4(n1018), .Z(n2204) );
  oan211d1 U12756 ( .C1(n1187), .C2(n1240), .B(n1275), .A(n1327), .ZN(n2203)
         );
  aoim31d1 U12757 ( .B1(n1234), .B2(n1335), .B3(n2204), .A(n2203), .ZN(N10566)
         );
  nd02d0 U12758 ( .A1(n1309), .A2(num_images[6]), .ZN(n2207) );
  oai211d1 U12759 ( .C1(n959), .C2(n999), .A(n1066), .B(n1096), .ZN(n2206) );
  aoi31d1 U12760 ( .B1(n1154), .B2(n1290), .B3(n1192), .A(n1521), .ZN(n2205)
         );
  aon211d1 U12761 ( .C1(n2207), .C2(n2206), .B(n2205), .A(n1362), .ZN(N10551)
         );
  nr02d0 U12762 ( .A1(n1337), .A2(n1250), .ZN(n2209) );
  nd04d0 U12763 ( .A1(n1207), .A2(n1157), .A3(n1105), .A4(n1071), .ZN(n2208)
         );
  aoim22d1 U12764 ( .A1(n2209), .A2(n2208), .B1(n1336), .B2(n1291), .Z(N10536)
         );
  nd02d0 U12765 ( .A1(n1253), .A2(n1304), .ZN(n2212) );
  nd03d0 U12766 ( .A1(n1206), .A2(num_images[4]), .A3(n1285), .ZN(n2211) );
  aoi321d1 U12767 ( .C1(n974), .C2(n1091), .C3(n1000), .B1(n1108), .B2(n1053), 
        .A(n1590), .ZN(n2210) );
  aon211d1 U12768 ( .C1(n2212), .C2(n2211), .B(n2210), .A(n1362), .ZN(N10521)
         );
  ora211d1 U12769 ( .C1(n1002), .C2(n1059), .A(n1116), .B(n1155), .Z(n2214) );
  oan211d1 U12770 ( .C1(n1187), .C2(n1240), .B(n1275), .A(n1327), .ZN(n2213)
         );
  aoim31d1 U12771 ( .B1(n1231), .B2(n1324), .B3(n2214), .A(n2213), .ZN(N10506)
         );
  an02d0 U12772 ( .A1(n1114), .A2(n1069), .Z(n2215) );
  oan211d1 U12773 ( .C1(n967), .C2(n1004), .B(n1094), .A(n2215), .ZN(n2218) );
  nd02d0 U12774 ( .A1(n1253), .A2(n1304), .ZN(n2217) );
  aoi31d1 U12775 ( .B1(n1197), .B2(n1149), .B3(n1286), .A(n1580), .ZN(n2216)
         );
  aon211d1 U12776 ( .C1(n2218), .C2(n2217), .B(n2216), .A(n1362), .ZN(N10491)
         );
  aoi311d1 U12777 ( .C1(n1158), .C2(n1095), .C3(n1195), .A(n1325), .B(n1225), 
        .ZN(n2219) );
  aoim21d1 U12778 ( .B1(n1299), .B2(n1344), .A(n2219), .ZN(N10476) );
  aoi31d1 U12779 ( .B1(n1018), .B2(n975), .B3(n1063), .A(n1110), .ZN(n2222) );
  nd02d0 U12780 ( .A1(n1253), .A2(n1305), .ZN(n2221) );
  aoi31d1 U12781 ( .B1(n1197), .B2(n1149), .B3(n1286), .A(n1590), .ZN(n2220)
         );
  aon211d1 U12782 ( .C1(n2222), .C2(n2221), .B(n2220), .A(n1362), .ZN(N10461)
         );
  an02d0 U12783 ( .A1(n1055), .A2(n1019), .Z(n2223) );
  aor22d1 U12784 ( .A1(n2223), .A2(n1147), .B1(n1111), .B2(n1154), .Z(n2225)
         );
  oan211d1 U12785 ( .C1(n1186), .C2(n1241), .B(n1275), .A(n1327), .ZN(n2224)
         );
  aoim31d1 U12786 ( .B1(n1250), .B2(n1329), .B3(n2225), .A(n2224), .ZN(N10446)
         );
  oan211d1 U12787 ( .C1(n966), .C2(n1004), .B(n1055), .A(n1098), .ZN(n2228) );
  nd02d0 U12788 ( .A1(n1252), .A2(n1304), .ZN(n2227) );
  aoi31d1 U12789 ( .B1(n1197), .B2(n1149), .B3(n1286), .A(n1580), .ZN(n2226)
         );
  aon211d1 U12790 ( .C1(n2228), .C2(n2227), .B(n2226), .A(n1362), .ZN(N10431)
         );
  nr02d0 U12791 ( .A1(n1336), .A2(n1249), .ZN(n2230) );
  oai211d1 U12792 ( .C1(n1042), .C2(n1091), .A(n1153), .B(n1189), .ZN(n2229)
         );
  aoim22d1 U12793 ( .A1(n2230), .A2(n2229), .B1(n1336), .B2(n1291), .Z(N10416)
         );
  an02d0 U12794 ( .A1(n1298), .A2(n1242), .Z(n2231) );
  aoi21d1 U12795 ( .B1(n1011), .B2(n964), .A(n2231), .ZN(n2234) );
  nr02d0 U12796 ( .A1(n1095), .A2(n1078), .ZN(n2233) );
  aoi31d1 U12797 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n2231), .ZN(n2232)
         );
  aon211d1 U12798 ( .C1(n2234), .C2(n2233), .B(n2232), .A(n1363), .ZN(N10401)
         );
  or02d0 U12799 ( .A1(n1027), .A2(n1037), .Z(n2235) );
  aor22d1 U12800 ( .A1(n1152), .A2(n2235), .B1(n1111), .B2(n1134), .Z(n2237)
         );
  oan211d1 U12801 ( .C1(n1187), .C2(n1242), .B(n1275), .A(n1327), .ZN(n2236)
         );
  aoim31d1 U12802 ( .B1(n1233), .B2(n1340), .B3(n2237), .A(n2236), .ZN(N10386)
         );
  an02d0 U12803 ( .A1(n1298), .A2(n1242), .Z(n2238) );
  nr02d0 U12804 ( .A1(n982), .A2(n2238), .ZN(n2241) );
  nr03d0 U12805 ( .A1(n1022), .A2(n1119), .A3(n1082), .ZN(n2240) );
  aoi31d1 U12806 ( .B1(n1154), .B2(n1290), .B3(n1193), .A(n2238), .ZN(n2239)
         );
  aon211d1 U12807 ( .C1(n2241), .C2(n2240), .B(n2239), .A(n1362), .ZN(N10371)
         );
  aoi321d1 U12808 ( .C1(n1145), .C2(n1272), .C3(n1181), .B1(n1277), .B2(n1229), 
        .A(n1337), .ZN(n2242) );
  nd03d0 U12809 ( .A1(n1180), .A2(n1140), .A3(n1301), .ZN(n2243) );
  oaim21d1 U12810 ( .B1(n1245), .B2(n1287), .A(n2243), .ZN(n2244) );
  nd04d0 U12811 ( .A1(n1091), .A2(n1073), .A3(n1025), .A4(n980), .ZN(n2246) );
  aoi21d1 U12812 ( .B1(n1278), .B2(n1189), .A(n2244), .ZN(n2245) );
  aon211d1 U12813 ( .C1(n2247), .C2(n2246), .B(n2245), .A(n1363), .ZN(N10341)
         );
  aor31d1 U12814 ( .B1(n1069), .B2(n1016), .B3(n1093), .A(n1147), .Z(n2249) );
  oan211d1 U12815 ( .C1(n1187), .C2(n1249), .B(n1275), .A(n1327), .ZN(n2248)
         );
  aoim31d1 U12816 ( .B1(n1234), .B2(n1347), .B3(n2249), .A(n2248), .ZN(N10326)
         );
  nd03d0 U12817 ( .A1(n1203), .A2(n1134), .A3(n1281), .ZN(n2250) );
  oaim21d1 U12818 ( .B1(n1245), .B2(n1288), .A(n2250), .ZN(n2251) );
  oai211d1 U12819 ( .C1(n959), .C2(n1022), .A(n1066), .B(n1096), .ZN(n2253) );
  aoi21d1 U12820 ( .B1(n1278), .B2(n1192), .A(n2251), .ZN(n2252) );
  aon211d1 U12821 ( .C1(n2254), .C2(n2253), .B(n2252), .A(n1362), .ZN(N10311)
         );
  or02d0 U12822 ( .A1(n1334), .A2(n1248), .Z(n2255) );
  aoi321d1 U12823 ( .C1(n1102), .C2(n1047), .C3(n1208), .B1(n1148), .B2(n1188), 
        .A(n2255), .ZN(n2256) );
  aoim21d1 U12824 ( .B1(n1346), .B2(n1291), .A(n2256), .ZN(N10296) );
  nd03d0 U12825 ( .A1(n1186), .A2(n1151), .A3(n1280), .ZN(n2257) );
  oaim21d1 U12826 ( .B1(n1245), .B2(n1287), .A(n2257), .ZN(n2259) );
  aoi321d1 U12827 ( .C1(n974), .C2(n1091), .C3(n1017), .B1(n1107), .B2(n1053), 
        .A(n2259), .ZN(n2258) );
  aon211d1 U12828 ( .C1(n1181), .C2(n1295), .B(n2259), .A(n2261), .ZN(n2260)
         );
  nd12d0 U12829 ( .A1(n1350), .A2(n2260), .ZN(N10281) );
  oan211d1 U12830 ( .C1(n1186), .C2(n1254), .B(n1275), .A(n1327), .ZN(n2262)
         );
  aoim31d1 U12831 ( .B1(n1234), .B2(n1338), .B3(n1865), .A(n2262), .ZN(N10266)
         );
  nd03d0 U12832 ( .A1(n1202), .A2(n1156), .A3(n1288), .ZN(n2263) );
  oaim21d1 U12833 ( .B1(n1245), .B2(n1288), .A(n2263), .ZN(n2266) );
  oai21d1 U12834 ( .B1(n974), .B2(n1009), .A(n1105), .ZN(n2264) );
  oaim2m11d1 U12835 ( .C1(n1114), .C2(n1064), .B(n2266), .A(n2264), .ZN(n2265)
         );
  aon211d1 U12836 ( .C1(n1180), .C2(n1282), .B(n2266), .A(n2265), .ZN(n2267)
         );
  nd12d0 U12837 ( .A1(n1350), .A2(n2267), .ZN(N10251) );
  nr02d0 U12838 ( .A1(n1331), .A2(n1249), .ZN(n2269) );
  oai21d1 U12839 ( .B1(n1101), .B2(n1139), .A(n1206), .ZN(n2268) );
  aoim22d1 U12840 ( .A1(n2269), .A2(n2268), .B1(n1294), .B2(n1332), .Z(N10236)
         );
  nd03d0 U12841 ( .A1(n1195), .A2(n1155), .A3(n1298), .ZN(n2270) );
  oaim21d1 U12842 ( .B1(n1244), .B2(n1287), .A(n2270), .ZN(n2272) );
  aor311d1 U12843 ( .C1(n1017), .C2(n975), .C3(n1051), .A(n2272), .B(n1116), 
        .Z(n2271) );
  aon211d1 U12844 ( .C1(n1181), .C2(n1303), .B(n2272), .A(n2271), .ZN(n2273)
         );
  nd12d0 U12845 ( .A1(n1350), .A2(n2273), .ZN(N10221) );
  aoi21d1 U12846 ( .B1(n1058), .B2(n1006), .A(n1110), .ZN(n2276) );
  nr03d0 U12847 ( .A1(num_images[4]), .A2(n1347), .A3(n1242), .ZN(n2275) );
  oai21d1 U12848 ( .B1(n1200), .B2(n1231), .A(n1281), .ZN(n2274) );
  aoi22d1 U12849 ( .A1(n2276), .A2(n2275), .B1(n2274), .B2(n1357), .ZN(N10206)
         );
  oan211d1 U12850 ( .C1(n967), .C2(n1003), .B(n1055), .A(n1099), .ZN(n2280) );
  nd03d0 U12851 ( .A1(n1183), .A2(n1159), .A3(n1278), .ZN(n2277) );
  oaim21d1 U12852 ( .B1(n1245), .B2(n1287), .A(n2277), .ZN(n2278) );
  aoi21d1 U12853 ( .B1(n1279), .B2(n1193), .A(n2278), .ZN(n2279) );
  aon211d1 U12854 ( .C1(n2280), .C2(n2281), .B(n2279), .A(n1362), .ZN(N10191)
         );
  or02d0 U12855 ( .A1(n1079), .A2(n1117), .Z(n2282) );
  aoi22d1 U12856 ( .A1(n1181), .A2(n2282), .B1(n1144), .B2(n1177), .ZN(n2284)
         );
  nr02d0 U12857 ( .A1(n1325), .A2(n1249), .ZN(n2283) );
  aoim22d1 U12858 ( .A1(n2284), .A2(n2283), .B1(n1336), .B2(n1291), .Z(N10176)
         );
  nd03d0 U12859 ( .A1(n1204), .A2(n1152), .A3(n1280), .ZN(n2285) );
  oaim21d1 U12860 ( .B1(n1245), .B2(n1287), .A(n2285), .ZN(n2288) );
  or02d0 U12861 ( .A1(n1120), .A2(n1086), .Z(n2286) );
  aor211d1 U12862 ( .C1(n1016), .C2(n965), .A(n2286), .B(n2288), .Z(n2287) );
  aon211d1 U12863 ( .C1(n1180), .C2(n1274), .B(n2288), .A(n2287), .ZN(n2289)
         );
  nd12d0 U12864 ( .A1(n1350), .A2(n2289), .ZN(N10161) );
  nr03d0 U12865 ( .A1(n1022), .A2(n1119), .A3(n1077), .ZN(n2292) );
  nr03d0 U12866 ( .A1(n1148), .A2(n1347), .A3(n1256), .ZN(n2291) );
  oai21d1 U12867 ( .B1(n1191), .B2(n1231), .A(n1281), .ZN(n2290) );
  aoi22d1 U12868 ( .A1(n2292), .A2(n2291), .B1(n2290), .B2(n1357), .ZN(N10146)
         );
  nd03d0 U12869 ( .A1(n1205), .A2(n1138), .A3(n1282), .ZN(n2293) );
  oaim21d1 U12870 ( .B1(n1244), .B2(n1287), .A(n2293), .ZN(n2296) );
  or02d0 U12871 ( .A1(n1093), .A2(n1082), .Z(n2294) );
  or04d0 U12872 ( .A1(n1021), .A2(n2294), .A3(n977), .A4(n2296), .Z(n2295) );
  aon211d1 U12873 ( .C1(n1181), .C2(n1301), .B(n2296), .A(n2295), .ZN(n2297)
         );
  nd12d0 U12874 ( .A1(n1350), .A2(n2297), .ZN(N10131) );
  oan211d1 U12875 ( .C1(n1228), .C2(n1181), .B(n1275), .A(n1326), .ZN(n2298)
         );
  aoi22d1 U12876 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1178), .ZN(n2301)
         );
  nd04d0 U12877 ( .A1(num_images[3]), .A2(n1073), .A3(n1024), .A4(n980), .ZN(
        n2300) );
  aoi21d1 U12878 ( .B1(n1143), .B2(n1298), .A(n1677), .ZN(n2299) );
  aon211d1 U12879 ( .C1(n2301), .C2(n2300), .B(n2299), .A(n1363), .ZN(N10101)
         );
  an04d0 U12880 ( .A1(n1158), .A2(n1114), .A3(n1074), .A4(n1019), .Z(n2302) );
  nr04d0 U12881 ( .A1(n1341), .A2(n1252), .A3(n1182), .A4(n2302), .ZN(n2303)
         );
  aoim21d1 U12882 ( .B1(n1300), .B2(n1333), .A(n2303), .ZN(N10086) );
  aoi22d1 U12883 ( .A1(n1226), .A2(n1272), .B1(n1285), .B2(n1178), .ZN(n2306)
         );
  oai211d1 U12884 ( .C1(n959), .C2(n999), .A(n1066), .B(n1096), .ZN(n2305) );
  aoi21d1 U12885 ( .B1(n1141), .B2(n1273), .A(n1677), .ZN(n2304) );
  aon211d1 U12886 ( .C1(n2306), .C2(n2305), .B(n2304), .A(n1363), .ZN(N10071)
         );
  aoi31d1 U12887 ( .B1(n1095), .B2(n1063), .B3(n1148), .A(n1204), .ZN(n2308)
         );
  nr02d0 U12888 ( .A1(n1337), .A2(n1250), .ZN(n2307) );
  aoim22d1 U12889 ( .A1(n2308), .A2(n2307), .B1(n1336), .B2(n1291), .Z(N10056)
         );
  aor22d1 U12890 ( .A1(n1237), .A2(n1282), .B1(n1292), .B2(n1207), .Z(n2309)
         );
  aoi321d1 U12891 ( .C1(n972), .C2(n1091), .C3(n1019), .B1(n1108), .B2(n1054), 
        .A(n2309), .ZN(n2311) );
  aoi21d1 U12892 ( .B1(n1141), .B2(n1273), .A(n2309), .ZN(n2310) );
  oai21d1 U12893 ( .B1(n2311), .B2(n2310), .A(n1361), .ZN(N10041) );
  ora211d1 U12894 ( .C1(n1002), .C2(n1059), .A(n1116), .B(n1155), .Z(n2312) );
  nr04d0 U12895 ( .A1(n1341), .A2(n1252), .A3(num_images[5]), .A4(n2312), .ZN(
        n2313) );
  aoim21d1 U12896 ( .B1(n1309), .B2(n1345), .A(n2313), .ZN(N10026) );
  aoi22d1 U12897 ( .A1(n1225), .A2(n1272), .B1(n1285), .B2(n1178), .ZN(n2314)
         );
  oai21d1 U12898 ( .B1(n974), .B2(n1009), .A(n1105), .ZN(n2315) );
  oaim211d1 U12899 ( .C1(n1113), .C2(n1067), .A(n2315), .B(n2314), .ZN(n2316)
         );
  aon211d1 U12900 ( .C1(n1138), .C2(n1278), .B(n1677), .A(n2316), .ZN(n2317)
         );
  nd12d0 U12901 ( .A1(n1350), .A2(n2317), .ZN(N10011) );
  aoi21d1 U12902 ( .B1(n1141), .B2(n1113), .A(n1178), .ZN(n2319) );
  nr02d0 U12903 ( .A1(n1325), .A2(n1249), .ZN(n2318) );
  aoim22d1 U12904 ( .A1(n2319), .A2(n2318), .B1(n1293), .B2(n1332), .Z(N9996)
         );
  aor22d1 U12905 ( .A1(n1238), .A2(n1283), .B1(n1292), .B2(n1197), .Z(n2321)
         );
  aor311d1 U12906 ( .C1(n1017), .C2(n976), .C3(n1050), .A(n1104), .B(n2321), 
        .Z(n2320) );
  aon211d1 U12907 ( .C1(n1149), .C2(n1302), .B(n2321), .A(n2320), .ZN(n2322)
         );
  nd12d0 U12908 ( .A1(n1350), .A2(n2322), .ZN(N9981) );
  or03d0 U12909 ( .A1(n1348), .A2(n1239), .A3(n1190), .Z(n2323) );
  aoi321d1 U12910 ( .C1(n1059), .C2(n1002), .C3(n1134), .B1(n1107), .B2(n1136), 
        .A(n2323), .ZN(n2324) );
  aoim21d1 U12911 ( .B1(n1296), .B2(n1329), .A(n2324), .ZN(N9966) );
  oan211d1 U12912 ( .C1(n967), .C2(n1005), .B(n1056), .A(n1098), .ZN(n2327) );
  aoi22d1 U12913 ( .A1(n1226), .A2(n1272), .B1(n1284), .B2(n1177), .ZN(n2326)
         );
  aoi21d1 U12914 ( .B1(n1142), .B2(n1273), .A(n2328), .ZN(n2325) );
  aon211d1 U12915 ( .C1(n2327), .C2(n2326), .B(n2325), .A(n1363), .ZN(N9951)
         );
  oan211d1 U12916 ( .C1(n1052), .C2(n1094), .B(n1137), .A(n1189), .ZN(n2330)
         );
  nr02d0 U12917 ( .A1(n1335), .A2(n1250), .ZN(n2329) );
  aoim22d1 U12918 ( .A1(n2330), .A2(n2329), .B1(n1336), .B2(n1291), .Z(N9936)
         );
  aor22d1 U12919 ( .A1(n1237), .A2(n1283), .B1(n1292), .B2(n1201), .Z(n2331)
         );
  aoi21d1 U12920 ( .B1(n1011), .B2(n964), .A(n2331), .ZN(n2334) );
  nr02d0 U12921 ( .A1(n1113), .A2(n1079), .ZN(n2333) );
  aoi21d1 U12922 ( .B1(n1142), .B2(n1276), .A(n2331), .ZN(n2332) );
  aon211d1 U12923 ( .C1(n2334), .C2(n2333), .B(n2332), .A(n1363), .ZN(N9921)
         );
  or02d0 U12924 ( .A1(n1027), .A2(n1039), .Z(n2335) );
  aoi22d1 U12925 ( .A1(n1132), .A2(n2335), .B1(n1106), .B2(n1134), .ZN(n2337)
         );
  nr03d0 U12926 ( .A1(n1203), .A2(n1347), .A3(n1256), .ZN(n2336) );
  aoim22d1 U12927 ( .A1(n2337), .A2(n2336), .B1(n1293), .B2(n1333), .Z(N9906)
         );
  aor22d1 U12928 ( .A1(n1237), .A2(n1283), .B1(n1292), .B2(n1182), .Z(n2338)
         );
  nr02d0 U12929 ( .A1(n982), .A2(n2338), .ZN(n2341) );
  nr03d0 U12930 ( .A1(n1021), .A2(n1119), .A3(n1078), .ZN(n2340) );
  aoi21d1 U12931 ( .B1(n1142), .B2(n1284), .A(n2338), .ZN(n2339) );
  aon211d1 U12932 ( .C1(n2341), .C2(n2340), .B(n2339), .A(n1363), .ZN(N9891)
         );
  oan211d1 U12933 ( .C1(n1135), .C2(n1181), .B(n1275), .A(n1327), .ZN(n2342)
         );
  oaim21d1 U12934 ( .B1(n1245), .B2(n1287), .A(n2342), .ZN(N9876) );
  an04d0 U12935 ( .A1(n1098), .A2(n1042), .A3(n1020), .A4(n978), .Z(n2343) );
  or04d0 U12936 ( .A1(n1158), .A2(n2343), .A3(n1239), .A4(n1192), .Z(n2344) );
  aor21d1 U12937 ( .B1(n1295), .B2(n2344), .A(n1328), .Z(N9861) );
  aoi31d1 U12938 ( .B1(n1068), .B2(n1015), .B3(n1107), .A(n1149), .ZN(n2346)
         );
  nr03d0 U12939 ( .A1(n1204), .A2(n1348), .A3(n1256), .ZN(n2345) );
  aoim22d1 U12940 ( .A1(n2346), .A2(n2345), .B1(n1294), .B2(n1333), .Z(N9846)
         );
  ora211d1 U12941 ( .C1(n963), .C2(n1013), .A(n1052), .B(n1094), .Z(n2347) );
  or04d0 U12942 ( .A1(n1158), .A2(n2347), .A3(n1238), .A4(n1177), .Z(n2348) );
  aor21d1 U12943 ( .B1(n1295), .B2(n2348), .A(n1328), .Z(N9831) );
  aoi21d1 U12944 ( .B1(n1100), .B2(n1050), .A(n1144), .ZN(n2350) );
  nr03d0 U12945 ( .A1(n1204), .A2(n1348), .A3(n1256), .ZN(n2349) );
  aoim22d1 U12946 ( .A1(n2350), .A2(n2349), .B1(n1336), .B2(n1291), .Z(N9816)
         );
  nd03d0 U12947 ( .A1(n982), .A2(n1102), .A3(n1028), .ZN(n2352) );
  nr03d0 U12948 ( .A1(n1153), .A2(n1228), .A3(n1208), .ZN(n2351) );
  oaim211d1 U12949 ( .C1(n1114), .C2(n1067), .A(n2352), .B(n2351), .ZN(n2353)
         );
  aor21d1 U12950 ( .B1(n1295), .B2(n2353), .A(n1328), .Z(N9801) );
  oan211d1 U12951 ( .C1(n1006), .C2(n1047), .B(n1094), .A(n1140), .ZN(n2355)
         );
  nr03d0 U12952 ( .A1(n1203), .A2(n1347), .A3(n1256), .ZN(n2354) );
  aoim22d1 U12953 ( .A1(n2355), .A2(n2354), .B1(n1293), .B2(n1333), .Z(N9786)
         );
  oai21d1 U12954 ( .B1(n974), .B2(n1009), .A(n1104), .ZN(n2357) );
  nr03d0 U12955 ( .A1(n1151), .A2(n1232), .A3(n1208), .ZN(n2356) );
  oaim211d1 U12956 ( .C1(n1114), .C2(n1067), .A(n2357), .B(n2356), .ZN(n2358)
         );
  nr02d0 U12957 ( .A1(n1162), .A2(n1117), .ZN(n2360) );
  nr03d0 U12958 ( .A1(n1204), .A2(n1348), .A3(n1240), .ZN(n2359) );
  aoim22d1 U12959 ( .A1(n2360), .A2(n2359), .B1(n1293), .B2(n1333), .Z(N9756)
         );
  aoi31d1 U12960 ( .B1(n1018), .B2(n975), .B3(n1063), .A(n1110), .ZN(n2362) );
  nr03d0 U12961 ( .A1(n1142), .A2(n1253), .A3(n1198), .ZN(n2361) );
  aon211d1 U12962 ( .C1(n2362), .C2(n2361), .B(n1310), .A(n1363), .ZN(N9741)
         );
  aoi211d1 U12963 ( .C1(n1062), .C2(n1008), .A(n1145), .B(n1089), .ZN(n2364)
         );
  nr03d0 U12964 ( .A1(n1204), .A2(n1347), .A3(n1226), .ZN(n2363) );
  aoim22d1 U12965 ( .A1(n2364), .A2(n2363), .B1(n1293), .B2(n1332), .Z(N9726)
         );
  oan211d1 U12966 ( .C1(n967), .C2(n1005), .B(n1057), .A(n1097), .ZN(n2366) );
  nr03d0 U12967 ( .A1(n1160), .A2(n1252), .A3(n1208), .ZN(n2365) );
  aon211d1 U12968 ( .C1(n2366), .C2(n2365), .B(n1271), .A(n1363), .ZN(N9711)
         );
  nr03d0 U12969 ( .A1(n1074), .A2(n1145), .A3(n1112), .ZN(n2368) );
  nr03d0 U12970 ( .A1(n1203), .A2(n1347), .A3(n1239), .ZN(n2367) );
  aoim22d1 U12971 ( .A1(n2368), .A2(n2367), .B1(n1336), .B2(n1291), .Z(N9696)
         );
  aoi211d1 U12972 ( .C1(n1014), .C2(n968), .A(n1102), .B(n1045), .ZN(n2370) );
  nr03d0 U12973 ( .A1(n1143), .A2(num_images[6]), .A3(n1208), .ZN(n2369) );
  aon211d1 U12974 ( .C1(n2370), .C2(n2369), .B(n1323), .A(n1363), .ZN(N9681)
         );
  nr03d0 U12975 ( .A1(n1022), .A2(n1119), .A3(n1074), .ZN(n2372) );
  nr04d0 U12976 ( .A1(n1341), .A2(n1252), .A3(num_images[5]), .A4(n1161), .ZN(
        n2371) );
  aoim22d1 U12977 ( .A1(n2372), .A2(n2371), .B1(n1293), .B2(n1333), .Z(N9666)
         );
  nr03d0 U12978 ( .A1(n979), .A2(n1071), .A3(n1027), .ZN(n2374) );
  nr04d0 U12979 ( .A1(n1230), .A2(n1204), .A3(n1163), .A4(num_images[3]), .ZN(
        n2373) );
  aon211d1 U12980 ( .C1(n2374), .C2(n2373), .B(n1321), .A(n1363), .ZN(N9652)
         );
  or02d0 U12981 ( .A1(n1299), .A2(n1340), .Z(N9638) );
  nd04d0 U12982 ( .A1(n1112), .A2(n1073), .A3(n1024), .A4(n980), .ZN(n2376) );
  aoi31d1 U12983 ( .B1(n1195), .B2(n1150), .B3(n1236), .A(n1289), .ZN(n2375)
         );
  aon211d1 U12984 ( .C1(n2376), .C2(n1318), .B(n2375), .A(n1364), .ZN(N9624)
         );
  nr02d0 U12985 ( .A1(N11556), .A2(n1306), .ZN(n2379) );
  nd04d0 U12986 ( .A1(n1162), .A2(n1114), .A3(n1073), .A4(n1023), .ZN(n2378)
         );
  nd02d0 U12987 ( .A1(n1252), .A2(n1202), .ZN(n2377) );
  aoi22d1 U12988 ( .A1(n2379), .A2(n2378), .B1(n2379), .B2(n2377), .ZN(N9610)
         );
  oai211d1 U12989 ( .C1(n960), .C2(n999), .A(n1064), .B(n1096), .ZN(n2381) );
  aoi31d1 U12990 ( .B1(n1196), .B2(n1150), .B3(n1236), .A(n1287), .ZN(n2380)
         );
  aon211d1 U12991 ( .C1(n2381), .C2(n1320), .B(n2380), .A(n1363), .ZN(N9596)
         );
  an04d0 U12992 ( .A1(n1202), .A2(n1156), .A3(n1116), .A4(n1069), .Z(n2383) );
  nr03d0 U12993 ( .A1(n1250), .A2(n1347), .A3(num_images[7]), .ZN(n2382) );
  aoim31d1 U12994 ( .B1(n1282), .B2(n1348), .B3(n2383), .A(n2382), .ZN(N9582)
         );
  nd03d0 U12995 ( .A1(n1185), .A2(n1132), .A3(n1257), .ZN(n2385) );
  aoi321d1 U12996 ( .C1(n973), .C2(n1087), .C3(n1000), .B1(n1108), .B2(n1054), 
        .A(n1294), .ZN(n2384) );
  aon211d1 U12997 ( .C1(n2385), .C2(n1271), .B(n2384), .A(n1361), .ZN(N9568)
         );
  nr02d0 U12998 ( .A1(n1349), .A2(n1306), .ZN(n2388) );
  oai211d1 U12999 ( .C1(n998), .C2(n1043), .A(n1111), .B(n1140), .ZN(n2387) );
  nd02d0 U13000 ( .A1(n1252), .A2(n1202), .ZN(n2386) );
  aoi22d1 U13001 ( .A1(n2388), .A2(n2387), .B1(n2388), .B2(n2386), .ZN(N9554)
         );
  aoi21d1 U13002 ( .B1(n1100), .B2(n1049), .A(n1289), .ZN(n2391) );
  oai21d1 U13003 ( .B1(N6867), .B2(n1010), .A(n1104), .ZN(n2390) );
  aoi31d1 U13004 ( .B1(n1195), .B2(n1151), .B3(n1236), .A(n1289), .ZN(n2389)
         );
  aon211d1 U13005 ( .C1(n2391), .C2(n2390), .B(n2389), .A(n1364), .ZN(N9540)
         );
  an02d0 U13006 ( .A1(n1156), .A2(n1113), .Z(n2392) );
  aor311d1 U13007 ( .C1(n1239), .C2(n1194), .C3(n2392), .A(n1333), .B(n1279), 
        .Z(N9526) );
  nd03d0 U13008 ( .A1(num_images[5]), .A2(n1163), .A3(n1257), .ZN(n2394) );
  aoi311d1 U13009 ( .C1(n1001), .C2(n962), .C3(n1042), .A(n1274), .B(n1090), 
        .ZN(n2393) );
  aon211d1 U13010 ( .C1(n2394), .C2(n1318), .B(n2393), .A(n1364), .ZN(N9512)
         );
  nr02d0 U13011 ( .A1(n1338), .A2(n1307), .ZN(n2397) );
  nd02d0 U13012 ( .A1(n1252), .A2(n1202), .ZN(n2396) );
  aoi321d1 U13013 ( .C1(n1059), .C2(n1003), .C3(n1134), .B1(n1108), .B2(n1136), 
        .A(n2669), .ZN(n2395) );
  aoi21d1 U13014 ( .B1(n2397), .B2(n2396), .A(n2395), .ZN(N9498) );
  nr02d0 U13015 ( .A1(n1302), .A2(n1108), .ZN(n2400) );
  oai21d1 U13016 ( .B1(n974), .B2(n1010), .A(n1061), .ZN(n2399) );
  aoi31d1 U13017 ( .B1(n1195), .B2(n1151), .B3(n1235), .A(n1290), .ZN(n2398)
         );
  aon211d1 U13018 ( .C1(n2400), .C2(n2399), .B(n2398), .A(n1364), .ZN(N9484)
         );
  ora211d1 U13019 ( .C1(n1046), .C2(n1102), .A(n1157), .B(n1199), .Z(n2402) );
  nr03d0 U13020 ( .A1(n1251), .A2(n1348), .A3(n1284), .ZN(n2401) );
  aoim31d1 U13021 ( .B1(n1282), .B2(n1324), .B3(n2402), .A(n2401), .ZN(N9470)
         );
  aoi21d1 U13022 ( .B1(n1012), .B2(n964), .A(n1063), .ZN(n2405) );
  nr02d0 U13023 ( .A1(n1306), .A2(n1109), .ZN(n2404) );
  aoi31d1 U13024 ( .B1(n1196), .B2(n1150), .B3(n1235), .A(n1296), .ZN(n2403)
         );
  aon211d1 U13025 ( .C1(n2405), .C2(n2404), .B(n2403), .A(n1364), .ZN(N9456)
         );
  nd02d0 U13026 ( .A1(n1093), .A2(n1159), .ZN(n2409) );
  oai21d1 U13027 ( .B1(n1012), .B2(n1058), .A(n1146), .ZN(n2408) );
  nr02d0 U13028 ( .A1(n1342), .A2(n1306), .ZN(n2407) );
  aoi21d1 U13029 ( .B1(n1232), .B2(n1194), .A(n2539), .ZN(n2406) );
  aoi31d1 U13030 ( .B1(n2409), .B2(n2408), .B3(n2407), .A(n2406), .ZN(N9442)
         );
  nr02d0 U13031 ( .A1(n1026), .A2(n978), .ZN(n2412) );
  nr03d0 U13032 ( .A1(n1070), .A2(n1283), .A3(n1103), .ZN(n2411) );
  aoi31d1 U13033 ( .B1(n1195), .B2(n1150), .B3(n1236), .A(n1289), .ZN(n2410)
         );
  aon211d1 U13034 ( .C1(n2412), .C2(n2411), .B(n2410), .A(n1364), .ZN(N9428)
         );
  aor311d1 U13035 ( .C1(n1195), .C2(n1151), .C3(n1227), .A(n1336), .B(n1273), 
        .Z(N9414) );
  aoi31d1 U13036 ( .B1(n1195), .B2(n1150), .B3(n1235), .A(n1289), .ZN(n2415)
         );
  nd04d0 U13037 ( .A1(n1120), .A2(n1073), .A3(n1024), .A4(n980), .ZN(n2414) );
  aoi21d1 U13038 ( .B1(n1233), .B2(n1179), .A(n2433), .ZN(n2413) );
  aon211d1 U13039 ( .C1(n2415), .C2(n2414), .B(n2413), .A(n1364), .ZN(N9400)
         );
  aoi31d1 U13040 ( .B1(n1068), .B2(n1015), .B3(n1107), .A(n1149), .ZN(n2418)
         );
  nr02d0 U13041 ( .A1(n1326), .A2(n1306), .ZN(n2417) );
  nd02d0 U13042 ( .A1(n1253), .A2(n1202), .ZN(n2416) );
  aoi22d1 U13043 ( .A1(n2418), .A2(n2417), .B1(n2417), .B2(n2416), .ZN(N9386)
         );
  aoi31d1 U13044 ( .B1(n1195), .B2(n1149), .B3(n1236), .A(n1289), .ZN(n2421)
         );
  oai211d1 U13045 ( .C1(n960), .C2(n1019), .A(n1066), .B(n1096), .ZN(n2420) );
  aoi21d1 U13046 ( .B1(n1233), .B2(n1191), .A(n1755), .ZN(n2419) );
  aon211d1 U13047 ( .C1(n2421), .C2(n2420), .B(n2419), .A(n1364), .ZN(N9372)
         );
  or02d0 U13048 ( .A1(n1276), .A2(n1340), .Z(n2422) );
  aoi321d1 U13049 ( .C1(n1101), .C2(n1046), .C3(n1177), .B1(n1148), .B2(n1188), 
        .A(n2422), .ZN(n2423) );
  aoim31d1 U13050 ( .B1(n1329), .B2(n1307), .B3(n1238), .A(n2423), .ZN(N9358)
         );
  aor31d1 U13051 ( .B1(n1198), .B2(n1152), .B3(n1228), .A(n1283), .Z(n2425) );
  aoi321d1 U13052 ( .C1(n974), .C2(n1091), .C3(n1000), .B1(n1108), .B2(n1054), 
        .A(n2425), .ZN(n2424) );
  aon211d1 U13053 ( .C1(n1180), .C2(n1252), .B(n2425), .A(n2427), .ZN(n2426)
         );
  nd12d0 U13054 ( .A1(n1349), .A2(n2426), .ZN(N9344) );
  oan211d1 U13055 ( .C1(n1007), .C2(n1048), .B(n1094), .A(n1140), .ZN(n2430)
         );
  nr02d0 U13056 ( .A1(n1327), .A2(n1307), .ZN(n2429) );
  nd02d0 U13057 ( .A1(n1253), .A2(n1202), .ZN(n2428) );
  aoi22d1 U13058 ( .A1(n2430), .A2(n2429), .B1(n2429), .B2(n2428), .ZN(N9330)
         );
  aor31d1 U13059 ( .B1(n1198), .B2(n1152), .B3(n1228), .A(n1283), .Z(n2433) );
  oai21d1 U13060 ( .B1(n957), .B2(n1010), .A(n1103), .ZN(n2431) );
  oaim2m11d1 U13061 ( .C1(n1114), .C2(n1064), .B(n2433), .A(n2431), .ZN(n2432)
         );
  aon211d1 U13062 ( .C1(n1180), .C2(n1223), .B(n2433), .A(n2432), .ZN(n2434)
         );
  nd12d0 U13063 ( .A1(n1349), .A2(n2434), .ZN(N9316) );
  or02d0 U13064 ( .A1(n1111), .A2(n1157), .Z(n2435) );
  aor311d1 U13065 ( .C1(n1195), .C2(n2435), .C3(n1228), .A(n1331), .B(n1276), 
        .Z(N9302) );
  aor31d1 U13066 ( .B1(n1198), .B2(n1152), .B3(n1228), .A(n1283), .Z(n2437) );
  aor311d1 U13067 ( .C1(n1017), .C2(n976), .C3(n1051), .A(n2437), .B(n1099), 
        .Z(n2436) );
  aon211d1 U13068 ( .C1(n1181), .C2(n1223), .B(n2437), .A(n2436), .ZN(n2438)
         );
  nd12d0 U13069 ( .A1(n1349), .A2(n2438), .ZN(N9288) );
  nr02d0 U13070 ( .A1(n1342), .A2(n1307), .ZN(n2439) );
  oaim21d1 U13071 ( .B1(n1086), .B2(n1015), .A(n2439), .ZN(n2441) );
  aoi21d1 U13072 ( .B1(n1233), .B2(n1185), .A(n2580), .ZN(n2440) );
  aoim31d1 U13073 ( .B1(n1146), .B2(n1115), .B3(n2441), .A(n2440), .ZN(N9274)
         );
  oan211d1 U13074 ( .C1(n965), .C2(n1003), .B(n1055), .A(n1098), .ZN(n2444) );
  aoi31d1 U13075 ( .B1(n1196), .B2(n1151), .B3(n1232), .A(n1306), .ZN(n2443)
         );
  aoi21d1 U13076 ( .B1(n1233), .B2(n1185), .A(n1765), .ZN(n2442) );
  aon211d1 U13077 ( .C1(n2444), .C2(n2443), .B(n2442), .A(n1364), .ZN(N9260)
         );
  or02d0 U13078 ( .A1(n1076), .A2(n1117), .Z(n2445) );
  aor22d1 U13079 ( .A1(n1194), .A2(n2445), .B1(n1153), .B2(n1179), .Z(n2447)
         );
  nr03d0 U13080 ( .A1(n1251), .A2(n1347), .A3(num_images[7]), .ZN(n2446) );
  aoim31d1 U13081 ( .B1(n1282), .B2(n1324), .B3(n2447), .A(n2446), .ZN(N9246)
         );
  aor31d1 U13082 ( .B1(n1199), .B2(n1152), .B3(n1228), .A(n1283), .Z(n2450) );
  or02d0 U13083 ( .A1(n1094), .A2(n1078), .Z(n2448) );
  aor211d1 U13084 ( .C1(n1016), .C2(n964), .A(n2448), .B(n2450), .Z(n2449) );
  aon211d1 U13085 ( .C1(n1180), .C2(n1223), .B(n2450), .A(n2449), .ZN(n2451)
         );
  nd12d0 U13086 ( .A1(n1349), .A2(n2451), .ZN(N9232) );
  nr02d0 U13087 ( .A1(n1333), .A2(n1307), .ZN(n2454) );
  nr03d0 U13088 ( .A1(n1070), .A2(n1137), .A3(n1092), .ZN(n2453) );
  aoi21d1 U13089 ( .B1(n1233), .B2(n1184), .A(n2568), .ZN(n2452) );
  aoi31d1 U13090 ( .B1(n2454), .B2(n1035), .B3(n2453), .A(n2452), .ZN(N9218)
         );
  aor31d1 U13091 ( .B1(n1199), .B2(n1152), .B3(n1228), .A(n1283), .Z(n2457) );
  or02d0 U13092 ( .A1(n1093), .A2(n1041), .Z(n2455) );
  or04d0 U13093 ( .A1(n1021), .A2(n2455), .A3(n977), .A4(n2457), .Z(n2456) );
  aon211d1 U13094 ( .C1(n1181), .C2(n1223), .B(n2457), .A(n2456), .ZN(n2458)
         );
  nd12d0 U13095 ( .A1(n1349), .A2(n2458), .ZN(N9204) );
  aor211d1 U13096 ( .C1(n1239), .C2(n1186), .A(n1348), .B(n1277), .Z(N9190) );
  aoi21d1 U13097 ( .B1(n1232), .B2(n1184), .A(n1299), .ZN(n2461) );
  nd04d0 U13098 ( .A1(n1120), .A2(n1072), .A3(n1024), .A4(n980), .ZN(n2460) );
  aoi21d1 U13099 ( .B1(n1143), .B2(n1221), .A(n2470), .ZN(n2459) );
  aon211d1 U13100 ( .C1(n2461), .C2(n2460), .B(n2459), .A(n1364), .ZN(N9176)
         );
  an02d0 U13101 ( .A1(n1069), .A2(n1019), .Z(n2462) );
  aoi31d1 U13102 ( .B1(n1154), .B2(n1110), .B3(n2462), .A(n1197), .ZN(n2464)
         );
  nr02d0 U13103 ( .A1(n1326), .A2(n1305), .ZN(n2463) );
  aoi22d1 U13104 ( .A1(n2464), .A2(n2463), .B1(n1222), .B2(n2463), .ZN(N9162)
         );
  aoi21d1 U13105 ( .B1(n1233), .B2(n1185), .A(n1308), .ZN(n2467) );
  oai211d1 U13106 ( .C1(n960), .C2(n1007), .A(n1066), .B(n1095), .ZN(n2466) );
  aoi21d1 U13107 ( .B1(n1142), .B2(num_images[6]), .A(n1829), .ZN(n2465) );
  aon211d1 U13108 ( .C1(n2467), .C2(n2466), .B(n2465), .A(n1364), .ZN(N9148)
         );
  aor31d1 U13109 ( .B1(n1112), .B2(n1064), .B3(n1136), .A(n1199), .Z(n2469) );
  nr03d0 U13110 ( .A1(n1251), .A2(n1347), .A3(n1270), .ZN(n2468) );
  aoim31d1 U13111 ( .B1(n1281), .B2(n1324), .B3(n2469), .A(n2468), .ZN(N9134)
         );
  aor21d1 U13112 ( .B1(n1241), .B2(n1191), .A(n1280), .Z(n2470) );
  aoi321d1 U13113 ( .C1(n974), .C2(n1090), .C3(n1000), .B1(n1109), .B2(n1053), 
        .A(n2470), .ZN(n2472) );
  aoi21d1 U13114 ( .B1(n1143), .B2(n1245), .A(n2470), .ZN(n2471) );
  oai21d1 U13115 ( .B1(n2472), .B2(n2471), .A(n1361), .ZN(N9120) );
  or02d0 U13116 ( .A1(n1027), .A2(n1075), .Z(n2473) );
  aoi31d1 U13117 ( .B1(n1096), .B2(n2473), .B3(n1148), .A(n1199), .ZN(n2475)
         );
  nr02d0 U13118 ( .A1(n1324), .A2(n1305), .ZN(n2474) );
  aoi22d1 U13119 ( .A1(n2475), .A2(n2474), .B1(n1269), .B2(n2474), .ZN(N9106)
         );
  aoi21d1 U13120 ( .B1(n1232), .B2(n1185), .A(n1290), .ZN(n2476) );
  oai21d1 U13121 ( .B1(n974), .B2(n1011), .A(n1103), .ZN(n2477) );
  oaim211d1 U13122 ( .C1(n1113), .C2(n1068), .A(n2477), .B(n2476), .ZN(n2478)
         );
  aon211d1 U13123 ( .C1(n1140), .C2(n1223), .B(n2499), .A(n2478), .ZN(n2479)
         );
  nd12d0 U13124 ( .A1(n1349), .A2(n2479), .ZN(N9092) );
  nd03d0 U13125 ( .A1(n1112), .A2(n1256), .A3(n1158), .ZN(n2481) );
  nr02d0 U13126 ( .A1(n1334), .A2(n1305), .ZN(n2480) );
  oaim211d1 U13127 ( .C1(n1243), .C2(n1195), .A(n2481), .B(n2480), .ZN(N9078)
         );
  aor21d1 U13128 ( .B1(n1230), .B2(n1191), .A(n1280), .Z(n2483) );
  aor311d1 U13129 ( .C1(n1017), .C2(n976), .C3(n1051), .A(n1102), .B(n2483), 
        .Z(n2482) );
  aon211d1 U13130 ( .C1(n1152), .C2(n1223), .B(n2483), .A(n2482), .ZN(n2484)
         );
  nd12d0 U13131 ( .A1(n1349), .A2(n2484), .ZN(N9064) );
  or02d0 U13132 ( .A1(n1333), .A2(n1302), .Z(n2485) );
  aoi21d1 U13133 ( .B1(n1100), .B2(n1141), .A(n2485), .ZN(n2487) );
  aoi31d1 U13134 ( .B1(n1068), .B2(n1015), .B3(n1148), .A(n1191), .ZN(n2486)
         );
  aoim22d1 U13135 ( .A1(n2487), .A2(n2486), .B1(n1240), .B2(n2485), .Z(N9050)
         );
  oan211d1 U13136 ( .C1(n965), .C2(n1003), .B(n1056), .A(n1098), .ZN(n2490) );
  aoi21d1 U13137 ( .B1(n1232), .B2(n1184), .A(n1290), .ZN(n2489) );
  aoi21d1 U13138 ( .B1(n1142), .B2(n1221), .A(n2483), .ZN(n2488) );
  aon211d1 U13139 ( .C1(n2490), .C2(n2489), .B(n2488), .A(n1365), .ZN(N9036)
         );
  nr03d0 U13140 ( .A1(n1252), .A2(n1348), .A3(n1296), .ZN(n2491) );
  aoim31d1 U13141 ( .B1(n1281), .B2(n1324), .B3(n1999), .A(n2491), .ZN(N9022)
         );
  aor21d1 U13142 ( .B1(n1241), .B2(n1191), .A(n1280), .Z(n2492) );
  aoi21d1 U13143 ( .B1(n1012), .B2(n964), .A(n2492), .ZN(n2495) );
  nr02d0 U13144 ( .A1(n1090), .A2(n1077), .ZN(n2494) );
  aoi21d1 U13145 ( .B1(n1141), .B2(n1257), .A(n2492), .ZN(n2493) );
  aon211d1 U13146 ( .C1(n2495), .C2(n2494), .B(n2493), .A(n1365), .ZN(N9008)
         );
  or02d0 U13147 ( .A1(n1341), .A2(n1302), .Z(n2496) );
  aoi21d1 U13148 ( .B1(n1100), .B2(n1137), .A(n2496), .ZN(n2498) );
  oan211d1 U13149 ( .C1(n1007), .C2(n1048), .B(n1137), .A(n1189), .ZN(n2497)
         );
  aoim22d1 U13150 ( .A1(n2498), .A2(n2497), .B1(n1240), .B2(n2496), .Z(N8994)
         );
  aor21d1 U13151 ( .B1(n1241), .B2(n1191), .A(n1280), .Z(n2499) );
  nr02d0 U13152 ( .A1(n982), .A2(n2499), .ZN(n2502) );
  nr03d0 U13153 ( .A1(n1021), .A2(n1119), .A3(n1040), .ZN(n2501) );
  aoi21d1 U13154 ( .B1(n1141), .B2(n1257), .A(n2499), .ZN(n2500) );
  aon211d1 U13155 ( .C1(n2502), .C2(n2501), .B(n2500), .A(n1365), .ZN(N8980)
         );
  or02d0 U13156 ( .A1(n1163), .A2(n1185), .Z(n2503) );
  oan211d1 U13157 ( .C1(n1147), .C2(n1182), .B(n1229), .A(n1277), .ZN(n2505)
         );
  nd04d0 U13158 ( .A1(n1120), .A2(n1072), .A3(n1024), .A4(n980), .ZN(n2504) );
  aoi22d1 U13159 ( .A1(n2505), .A2(n2504), .B1(n2505), .B2(n1222), .ZN(n2506)
         );
  or02d0 U13160 ( .A1(n1340), .A2(n2506), .Z(N8952) );
  or02d0 U13161 ( .A1(n1350), .A2(n1302), .Z(n2507) );
  aoi31d1 U13162 ( .B1(n1068), .B2(n1015), .B3(n1106), .A(n2507), .ZN(n2509)
         );
  nr02d0 U13163 ( .A1(n1198), .A2(n1159), .ZN(n2508) );
  aoim22d1 U13164 ( .A1(n2509), .A2(n2508), .B1(n1240), .B2(n2507), .Z(N8938)
         );
  oan211d1 U13165 ( .C1(n1146), .C2(n1181), .B(n1229), .A(n1277), .ZN(n2511)
         );
  oai211d1 U13166 ( .C1(n960), .C2(n999), .A(n1065), .B(n1095), .ZN(n2510) );
  aoi22d1 U13167 ( .A1(n2511), .A2(n2510), .B1(n2511), .B2(n1269), .ZN(n2512)
         );
  or02d0 U13168 ( .A1(n1350), .A2(n2512), .Z(N8924) );
  or03d0 U13169 ( .A1(n1348), .A2(n1303), .A3(n1181), .Z(n2513) );
  aoi211d1 U13170 ( .C1(n1106), .C2(n1056), .A(n2513), .B(num_images[4]), .ZN(
        n2514) );
  aoim31d1 U13171 ( .B1(n1330), .B2(n1289), .B3(n1224), .A(n2514), .ZN(N8910)
         );
  oan211d1 U13172 ( .C1(n1158), .C2(n1182), .B(n1230), .A(n1277), .ZN(n2516)
         );
  aoi321d1 U13173 ( .C1(n973), .C2(n1091), .C3(n1016), .B1(n1108), .B2(n1054), 
        .A(n1883), .ZN(n2515) );
  aon211d1 U13174 ( .C1(n2516), .C2(n1266), .B(n2515), .A(n1365), .ZN(N8896)
         );
  or02d0 U13175 ( .A1(n1339), .A2(n1303), .Z(n2517) );
  oan211d1 U13176 ( .C1(n1007), .C2(n1048), .B(n1093), .A(n2517), .ZN(n2519)
         );
  nr02d0 U13177 ( .A1(n1201), .A2(n1160), .ZN(n2518) );
  aoim22d1 U13178 ( .A1(n2519), .A2(n2518), .B1(n1240), .B2(n2517), .Z(N8882)
         );
  oan211d1 U13179 ( .C1(n1145), .C2(n1182), .B(n1230), .A(n1277), .ZN(n2521)
         );
  oai21d1 U13180 ( .B1(n973), .B2(n1010), .A(n1105), .ZN(n2520) );
  oaim211d1 U13181 ( .C1(n1113), .C2(n1068), .A(n2521), .B(n2520), .ZN(n2522)
         );
  oan211d1 U13182 ( .C1(n1883), .C2(n1239), .B(n2522), .A(n1328), .ZN(n2523)
         );
  oai21d1 U13183 ( .B1(n1102), .B2(n1139), .A(n1232), .ZN(n2525) );
  nr02d0 U13184 ( .A1(n1328), .A2(n1306), .ZN(n2524) );
  oaim211d1 U13185 ( .C1(n1243), .C2(n1195), .A(n2525), .B(n2524), .ZN(N8854)
         );
  aor311d1 U13186 ( .C1(n1017), .C2(n975), .C3(n1050), .A(n1883), .B(n1115), 
        .Z(n2526) );
  oan211d1 U13187 ( .C1(n2546), .C2(n1221), .B(n2526), .A(n1328), .ZN(n2527)
         );
  or02d0 U13188 ( .A1(n1327), .A2(n1303), .Z(n2528) );
  aoi21d1 U13189 ( .B1(n1059), .B2(n1005), .A(n2528), .ZN(n2530) );
  nr03d0 U13190 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n2529) );
  aoim22d1 U13191 ( .A1(n2530), .A2(n2529), .B1(n1240), .B2(n2528), .Z(N8826)
         );
  oan211d1 U13192 ( .C1(n965), .C2(n1004), .B(n1057), .A(n1099), .ZN(n2532) );
  oan211d1 U13193 ( .C1(n1154), .C2(n1183), .B(n1229), .A(n1277), .ZN(n2531)
         );
  aoi22d1 U13194 ( .A1(n2532), .A2(n2531), .B1(n2531), .B2(n1268), .ZN(n2533)
         );
  or02d0 U13195 ( .A1(n1325), .A2(n2533), .Z(N8812) );
  or03d0 U13196 ( .A1(n1348), .A2(n1303), .A3(n1195), .Z(n2534) );
  nr04d0 U13197 ( .A1(n2534), .A2(n1070), .A3(n1162), .A4(n1099), .ZN(n2535)
         );
  aoim31d1 U13198 ( .B1(n1329), .B2(n1305), .B3(n1226), .A(n2535), .ZN(N8798)
         );
  oan211d1 U13199 ( .C1(n1134), .C2(n1182), .B(n1230), .A(n1277), .ZN(n2538)
         );
  oaim21d1 U13200 ( .B1(n1019), .B2(N6867), .A(n2538), .ZN(n2536) );
  nr03d0 U13201 ( .A1(n2536), .A2(n1119), .A3(n1080), .ZN(n2537) );
  aon211d1 U13202 ( .C1(n2538), .C2(n1258), .B(n2537), .A(n1365), .ZN(N8784)
         );
  or02d0 U13203 ( .A1(n1324), .A2(n1303), .Z(n2539) );
  nr03d0 U13204 ( .A1(n2539), .A2(n1071), .A3(n1028), .ZN(n2541) );
  nr03d0 U13205 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n2540) );
  aoim22d1 U13206 ( .A1(n2541), .A2(n2540), .B1(n1240), .B2(n2539), .Z(N8770)
         );
  oan211d1 U13207 ( .C1(n1144), .C2(n1182), .B(n1230), .A(n1277), .ZN(n2542)
         );
  or02d0 U13208 ( .A1(n1103), .A2(n1079), .Z(n2543) );
  or04d0 U13209 ( .A1(n1021), .A2(n2543), .A3(n977), .A4(n2546), .Z(n2544) );
  oan211d1 U13210 ( .C1(n2546), .C2(n1249), .B(n2544), .A(n1327), .ZN(n2545)
         );
  or03d0 U13211 ( .A1(n1348), .A2(n1303), .A3(n1247), .Z(N8744) );
  nr02d0 U13212 ( .A1(n1255), .A2(n1306), .ZN(n2549) );
  nd04d0 U13213 ( .A1(n1120), .A2(n1041), .A3(n1025), .A4(n980), .ZN(n2548) );
  aoi21d1 U13214 ( .B1(n1190), .B2(num_images[4]), .A(n2578), .ZN(n2547) );
  aon211d1 U13215 ( .C1(n2549), .C2(n2548), .B(n2547), .A(n1365), .ZN(N8731)
         );
  nd04d0 U13216 ( .A1(n1147), .A2(n1103), .A3(n1082), .A4(n1023), .ZN(n2552)
         );
  nr02d0 U13217 ( .A1(n1348), .A2(n1305), .ZN(n2551) );
  nr13d1 U13218 ( .A1(n2551), .A2(n1234), .A3(n1184), .ZN(n2550) );
  aoi31d1 U13219 ( .B1(n2552), .B2(n1266), .B3(n2551), .A(n2550), .ZN(N8718)
         );
  nr02d0 U13220 ( .A1(n1254), .A2(n1305), .ZN(n2555) );
  oai211d1 U13221 ( .C1(n961), .C2(n1024), .A(n1065), .B(n1094), .ZN(n2554) );
  aoi21d1 U13222 ( .B1(n1190), .B2(num_images[4]), .A(n2556), .ZN(n2553) );
  aon211d1 U13223 ( .C1(n2555), .C2(n2554), .B(n2553), .A(n1365), .ZN(N8705)
         );
  an04d0 U13224 ( .A1(n1202), .A2(n1156), .A3(n1116), .A4(n1069), .Z(n2557) );
  or04d0 U13225 ( .A1(n1238), .A2(n2557), .A3(n1334), .A4(n1282), .Z(N8692) );
  nr02d0 U13226 ( .A1(n1255), .A2(n1305), .ZN(n2560) );
  nd02d0 U13227 ( .A1(n1205), .A2(n1159), .ZN(n2559) );
  aoi321d1 U13228 ( .C1(n973), .C2(num_images[3]), .C3(n1020), .B1(n1109), 
        .B2(n1055), .A(n2556), .ZN(n2558) );
  aon211d1 U13229 ( .C1(n2560), .C2(n2559), .B(n2558), .A(n1365), .ZN(N8679)
         );
  oai211d1 U13230 ( .C1(n998), .C2(n1043), .A(n1111), .B(n1140), .ZN(n2563) );
  nr02d0 U13231 ( .A1(n1330), .A2(n1305), .ZN(n2562) );
  nr13d1 U13232 ( .A1(n2562), .A2(n1238), .A3(n1182), .ZN(n2561) );
  aoi31d1 U13233 ( .B1(n2563), .B2(n1267), .B3(n2562), .A(n2561), .ZN(N8666)
         );
  nr02d0 U13234 ( .A1(n1254), .A2(n1305), .ZN(n2564) );
  oai21d1 U13235 ( .B1(n972), .B2(n1011), .A(n1105), .ZN(n2565) );
  oaim211d1 U13236 ( .C1(n1113), .C2(n1067), .A(n2565), .B(n2564), .ZN(n2566)
         );
  aon211d1 U13237 ( .C1(n1180), .C2(n1141), .B(n1901), .A(n2566), .ZN(n2567)
         );
  nd12d0 U13238 ( .A1(n1350), .A2(n2567), .ZN(N8653) );
  or02d0 U13239 ( .A1(n1325), .A2(n1302), .Z(n2568) );
  aor311d1 U13240 ( .C1(n1154), .C2(n1110), .C3(n1186), .A(n1232), .B(n2568), 
        .Z(N8640) );
  or02d0 U13241 ( .A1(n1241), .A2(n1302), .Z(n2570) );
  aor311d1 U13242 ( .C1(n1017), .C2(n975), .C3(n1050), .A(n1120), .B(n2570), 
        .Z(n2569) );
  aon211d1 U13243 ( .C1(n1180), .C2(n1138), .B(n2570), .A(n2569), .ZN(n2571)
         );
  nd12d0 U13244 ( .A1(n1350), .A2(n2571), .ZN(N8627) );
  or02d0 U13245 ( .A1(n1345), .A2(n1302), .Z(n2574) );
  aor31d1 U13246 ( .B1(n1069), .B2(n1015), .B3(n1136), .A(n1235), .Z(n2572) );
  aoi211d1 U13247 ( .C1(n1100), .C2(n1138), .A(n2572), .B(n2574), .ZN(n2573)
         );
  aoim31d1 U13248 ( .B1(n1234), .B2(n1183), .B3(n2574), .A(n2573), .ZN(N8614)
         );
  oan211d1 U13249 ( .C1(n966), .C2(n1003), .B(n1057), .A(n1098), .ZN(n2577) );
  nr02d0 U13250 ( .A1(n1255), .A2(n1306), .ZN(n2576) );
  aoi21d1 U13251 ( .B1(n1190), .B2(n1132), .A(n2578), .ZN(n2575) );
  aon211d1 U13252 ( .C1(n2577), .C2(n2576), .B(n2575), .A(n1365), .ZN(N8601)
         );
  ora211d1 U13253 ( .C1(n1046), .C2(n1102), .A(n1135), .B(n1199), .Z(n2579) );
  aor211d1 U13254 ( .C1(n1004), .C2(n965), .A(n1089), .B(n1046), .Z(n2581) );
  or02d0 U13255 ( .A1(n1343), .A2(n1302), .Z(n2580) );
  aor311d1 U13256 ( .C1(n1153), .C2(n2581), .C3(n1186), .A(n1241), .B(n2580), 
        .Z(N8575) );
  nr02d0 U13257 ( .A1(n1348), .A2(n1306), .ZN(n2582) );
  aoi21d1 U13258 ( .B1(n1101), .B2(num_images[4]), .A(n2604), .ZN(n2585) );
  oan211d1 U13259 ( .C1(n1006), .C2(n1048), .B(n1138), .A(n1232), .ZN(n2584)
         );
  nr02d0 U13260 ( .A1(n1255), .A2(n1202), .ZN(n2583) );
  aoi22d1 U13261 ( .A1(n2585), .A2(n2584), .B1(n2583), .B2(n2582), .ZN(N8562)
         );
  or04d0 U13262 ( .A1(n1020), .A2(n977), .A3(n1111), .A4(n1062), .Z(n2587) );
  or02d0 U13263 ( .A1(n1336), .A2(n1302), .Z(n2586) );
  aor311d1 U13264 ( .C1(n1153), .C2(n2587), .C3(n1186), .A(n1228), .B(n2586), 
        .Z(N8549) );
  an02d0 U13265 ( .A1(n1201), .A2(n1155), .Z(n2588) );
  or04d0 U13266 ( .A1(n1231), .A2(n2588), .A3(n1334), .A4(n1282), .Z(N8536) );
  aoi211d1 U13267 ( .C1(n1192), .C2(n1139), .A(n1280), .B(n1253), .ZN(n2590)
         );
  nd04d0 U13268 ( .A1(n1120), .A2(n1072), .A3(n1025), .A4(n981), .ZN(n2589) );
  aoi22d1 U13269 ( .A1(n2590), .A2(n2589), .B1(n2590), .B2(n1217), .ZN(n2591)
         );
  or02d0 U13270 ( .A1(n1328), .A2(n2591), .Z(N8523) );
  or02d0 U13271 ( .A1(n1335), .A2(n1302), .Z(n2594) );
  or02d0 U13272 ( .A1(n1256), .A2(n1158), .Z(n2592) );
  aoi311d1 U13273 ( .C1(n1046), .C2(n1006), .C3(n1105), .A(n2592), .B(n2594), 
        .ZN(n2593) );
  aoim31d1 U13274 ( .B1(n1247), .B2(n1183), .B3(n2594), .A(n2593), .ZN(N8510)
         );
  aoi211d1 U13275 ( .C1(n1192), .C2(n1137), .A(n1281), .B(n1237), .ZN(n2596)
         );
  oai211d1 U13276 ( .C1(n961), .C2(n999), .A(n1065), .B(n1095), .ZN(n2595) );
  aoi22d1 U13277 ( .A1(n2596), .A2(n2595), .B1(n2596), .B2(n1217), .ZN(n2597)
         );
  or02d0 U13278 ( .A1(n1327), .A2(n2597), .Z(N8497) );
  nd03d0 U13279 ( .A1(n1040), .A2(n1209), .A3(n1100), .ZN(n2599) );
  nr03d0 U13280 ( .A1(n1251), .A2(n1347), .A3(n1289), .ZN(n2598) );
  oaim211d1 U13281 ( .C1(n1188), .C2(n1153), .A(n2599), .B(n2598), .ZN(N8484)
         );
  aoi321d1 U13282 ( .C1(n973), .C2(num_images[3]), .C3(num_images[1]), .B1(
        n1109), .B2(n1053), .A(n13), .ZN(n2600) );
  oan211d1 U13283 ( .C1(n13), .C2(n1181), .B(n2602), .A(n1326), .ZN(n2601) );
  or02d0 U13284 ( .A1(N11556), .A2(n1301), .Z(n2604) );
  oan211d1 U13285 ( .C1(n1007), .C2(n1048), .B(n1094), .A(n2604), .ZN(n2603)
         );
  nr03d0 U13286 ( .A1(n2604), .A2(n1251), .A3(n1175), .ZN(n2605) );
  aoim31d1 U13287 ( .B1(n1147), .B2(num_images[6]), .B3(n2606), .A(n2605), 
        .ZN(N8458) );
  aoi211d1 U13288 ( .C1(n1192), .C2(n1137), .A(n1280), .B(n1245), .ZN(n2608)
         );
  oai21d1 U13289 ( .B1(n973), .B2(n1010), .A(n1104), .ZN(n2607) );
  oaim211d1 U13290 ( .C1(n1113), .C2(n1068), .A(n2608), .B(n2607), .ZN(n2609)
         );
  oan211d1 U13291 ( .C1(n1944), .C2(n1181), .B(n2609), .A(n1326), .ZN(n2610)
         );
  oan211d1 U13292 ( .C1(n1093), .C2(num_images[4]), .B(n1188), .A(n1232), .ZN(
        n2612) );
  nr02d0 U13293 ( .A1(N11556), .A2(n1306), .ZN(n2611) );
  nd02d0 U13294 ( .A1(n2612), .A2(n2611), .ZN(N8432) );
  aor211d1 U13295 ( .C1(n1195), .C2(n1148), .A(n1293), .B(n1224), .Z(n2614) );
  aor311d1 U13296 ( .C1(n1017), .C2(n976), .C3(n1051), .A(n2614), .B(n1097), 
        .Z(n2613) );
  oan211d1 U13297 ( .C1(n2614), .C2(n1181), .B(n2613), .A(n1326), .ZN(n2615)
         );
  nr02d0 U13298 ( .A1(n1329), .A2(n1306), .ZN(n2616) );
  oaim21d1 U13299 ( .B1(n1075), .B2(n1014), .A(n2616), .ZN(n2617) );
  nr04d0 U13300 ( .A1(n2617), .A2(n1109), .A3(n1255), .A4(n1153), .ZN(n2618)
         );
  aoim31d1 U13301 ( .B1(n1235), .B2(n1184), .B3(n2586), .A(n2618), .ZN(N8406)
         );
  oan211d1 U13302 ( .C1(n965), .C2(n1003), .B(n1055), .A(n1098), .ZN(n2620) );
  aoi211d1 U13303 ( .C1(n1192), .C2(n1137), .A(n1280), .B(n1252), .ZN(n2619)
         );
  aoi22d1 U13304 ( .A1(n2620), .A2(n2619), .B1(n2619), .B2(n1217), .ZN(n2621)
         );
  or02d0 U13305 ( .A1(n1326), .A2(n2621), .Z(N8393) );
  oai21d1 U13306 ( .B1(n1060), .B2(n1096), .A(n1201), .ZN(n2623) );
  nr03d0 U13307 ( .A1(n1251), .A2(n1347), .A3(n1292), .ZN(n2622) );
  oaim211d1 U13308 ( .C1(n1200), .C2(n1153), .A(n2623), .B(n2622), .ZN(N8380)
         );
  or02d0 U13309 ( .A1(n1110), .A2(n1074), .Z(n2624) );
  oan211d1 U13310 ( .C1(n12), .C2(n1183), .B(n5), .A(n1327), .ZN(n2625) );
  or02d0 U13311 ( .A1(n1331), .A2(n1302), .Z(n2628) );
  or03d0 U13312 ( .A1(n1237), .A2(n1158), .A3(n1116), .Z(n2626) );
  nr04d0 U13313 ( .A1(n2626), .A2(n2628), .A3(n1086), .A4(n1023), .ZN(n2627)
         );
  aoim31d1 U13314 ( .B1(n1244), .B2(n1184), .B3(n2628), .A(n2627), .ZN(N8354)
         );
  nr04d0 U13315 ( .A1(n1089), .A2(n1070), .A3(n1026), .A4(n979), .ZN(n2631) );
  nd02d0 U13316 ( .A1(n1205), .A2(n1159), .ZN(n2630) );
  nr03d0 U13317 ( .A1(n1251), .A2(n1347), .A3(n1295), .ZN(n2629) );
  oai211d1 U13318 ( .C1(n2631), .C2(n1217), .A(n2630), .B(n2629), .ZN(N8342)
         );
  or04d0 U13319 ( .A1(n1227), .A2(n1200), .A3(n1334), .A4(n1282), .Z(N8330) );
  nr03d0 U13320 ( .A1(n1307), .A2(n1253), .A3(n1197), .ZN(n2633) );
  nd04d0 U13321 ( .A1(n1120), .A2(n1075), .A3(n1026), .A4(n982), .ZN(n2632) );
  aoi22d1 U13322 ( .A1(n2633), .A2(n2632), .B1(n1164), .B2(n2633), .ZN(n2634)
         );
  or02d0 U13323 ( .A1(n1344), .A2(n2634), .Z(N8318) );
  nd04d0 U13324 ( .A1(n1162), .A2(n1105), .A3(n1040), .A4(n1023), .ZN(n2636)
         );
  nr03d0 U13325 ( .A1(n1251), .A2(n1347), .A3(num_images[7]), .ZN(n2635) );
  nd13d1 U13326 ( .A1(n1182), .A2(n2636), .A3(n2635), .ZN(N8306) );
  oai21d1 U13327 ( .B1(n1013), .B2(n968), .A(n1061), .ZN(n2639) );
  nd02d0 U13328 ( .A1(n1161), .A2(n1096), .ZN(n2638) );
  nr03d0 U13329 ( .A1(n1251), .A2(n1346), .A3(n1301), .ZN(n2637) );
  oai211d1 U13330 ( .C1(n2639), .C2(n2638), .A(n1220), .B(n2637), .ZN(N8294)
         );
  or03d0 U13331 ( .A1(n1348), .A2(n1304), .A3(n1247), .Z(n2640) );
  aor311d1 U13332 ( .C1(n1112), .C2(n1064), .C3(n1159), .A(n1206), .B(n2640), 
        .Z(N8282) );
  aoi321d1 U13333 ( .C1(n972), .C2(num_images[3]), .C3(n1000), .B1(n1107), 
        .B2(n1054), .A(n8), .ZN(n2641) );
  oan211d1 U13334 ( .C1(n8), .C2(n1132), .B(n2643), .A(n1327), .ZN(n2642) );
  oai211d1 U13335 ( .C1(n998), .C2(n1044), .A(n1111), .B(n1139), .ZN(n2645) );
  nr03d0 U13336 ( .A1(n1250), .A2(n1346), .A3(n1270), .ZN(n2644) );
  nd13d1 U13337 ( .A1(n1190), .A2(n2645), .A3(n2644), .ZN(N8258) );
  nr03d0 U13338 ( .A1(n1307), .A2(n1253), .A3(n1199), .ZN(n2646) );
  oai21d1 U13339 ( .B1(n972), .B2(n1011), .A(n1104), .ZN(n2647) );
  oaim211d1 U13340 ( .C1(n1113), .C2(n1067), .A(n2647), .B(n2646), .ZN(n2648)
         );
  oan211d1 U13341 ( .C1(n1136), .C2(n2026), .B(n2648), .A(n1326), .ZN(n2649)
         );
  aoi21d1 U13342 ( .B1(n1144), .B2(n1102), .A(n1203), .ZN(n2651) );
  nr03d0 U13343 ( .A1(n1250), .A2(n1346), .A3(num_images[7]), .ZN(n2650) );
  nd02d0 U13344 ( .A1(n2651), .A2(n2650), .ZN(N8234) );
  or03d0 U13345 ( .A1(n1285), .A2(n1255), .A3(n1182), .Z(n2653) );
  aor311d1 U13346 ( .C1(n1016), .C2(n976), .C3(n1051), .A(n1097), .B(n2653), 
        .Z(n2652) );
  oan211d1 U13347 ( .C1(n1136), .C2(n2653), .B(n2652), .A(n1327), .ZN(n2654)
         );
  aoi21d1 U13348 ( .B1(n1144), .B2(n1117), .A(n1196), .ZN(n2656) );
  nr03d0 U13349 ( .A1(n1251), .A2(n1346), .A3(n1293), .ZN(n2655) );
  oaim311d1 U13350 ( .C1(n1016), .C2(n1153), .C3(n1061), .A(n2656), .B(n2655), 
        .ZN(N8210) );
  oan211d1 U13351 ( .C1(n966), .C2(n1005), .B(n1057), .A(n1098), .ZN(n2658) );
  nr03d0 U13352 ( .A1(n1307), .A2(n1253), .A3(n1192), .ZN(n2657) );
  aoi22d1 U13353 ( .A1(n2658), .A2(n2657), .B1(n1171), .B2(n2657), .ZN(n2659)
         );
  or02d0 U13354 ( .A1(n1326), .A2(n2659), .Z(N8198) );
  oan211d1 U13355 ( .C1(n1052), .C2(num_images[3]), .B(n1139), .A(n1189), .ZN(
        n2661) );
  nr03d0 U13356 ( .A1(n1251), .A2(n1346), .A3(num_images[7]), .ZN(n2660) );
  nd02d0 U13357 ( .A1(n2661), .A2(n2660), .ZN(N8186) );
  aoi211d1 U13358 ( .C1(n1014), .C2(n968), .A(n1102), .B(n1045), .ZN(n2663) );
  nr03d0 U13359 ( .A1(n1250), .A2(n1346), .A3(n1297), .ZN(n2662) );
  oai211d1 U13360 ( .C1(n2663), .C2(n1133), .A(n1210), .B(n2662), .ZN(N8174)
         );
  nr02d0 U13361 ( .A1(n1026), .A2(n1038), .ZN(n2666) );
  aoi21d1 U13362 ( .B1(n1143), .B2(n1114), .A(n1198), .ZN(n2665) );
  nr03d0 U13363 ( .A1(n1251), .A2(n1346), .A3(n1282), .ZN(n2664) );
  oai211d1 U13364 ( .C1(n2666), .C2(n1172), .A(n2665), .B(n2664), .ZN(N8162)
         );
  nr04d0 U13365 ( .A1(n1117), .A2(n1070), .A3(n1027), .A4(n979), .ZN(n2668) );
  nr03d0 U13366 ( .A1(n1250), .A2(n1346), .A3(n1294), .ZN(n2667) );
  oai211d1 U13367 ( .C1(n2668), .C2(n1164), .A(n1176), .B(n2667), .ZN(N8151)
         );
  or02d0 U13368 ( .A1(n1328), .A2(n1302), .Z(n2669) );
  nr02d0 U13369 ( .A1(n1207), .A2(n1160), .ZN(n2672) );
  nd04d0 U13370 ( .A1(n1092), .A2(n1072), .A3(n1026), .A4(n982), .ZN(n2671) );
  nr03d0 U13371 ( .A1(n1250), .A2(n1346), .A3(n1298), .ZN(n2670) );
  nd03d0 U13372 ( .A1(n2672), .A2(n2671), .A3(n2670), .ZN(N8129) );
  aor311d1 U13373 ( .C1(n1068), .C2(n1015), .C3(n1092), .A(n1196), .B(n1134), 
        .Z(n2673) );
  nr02d0 U13374 ( .A1(n1207), .A2(n1160), .ZN(n2676) );
  oai211d1 U13375 ( .C1(n998), .C2(n961), .A(n1065), .B(n1096), .ZN(n2675) );
  nr03d0 U13376 ( .A1(n1251), .A2(n1346), .A3(num_images[7]), .ZN(n2674) );
  nd03d0 U13377 ( .A1(n2676), .A2(n2675), .A3(n2674), .ZN(N8107) );
  aoi211d1 U13378 ( .C1(n1106), .C2(n1056), .A(n1192), .B(n1163), .ZN(n2678)
         );
  nr03d0 U13379 ( .A1(n1250), .A2(n1346), .A3(num_images[7]), .ZN(n2677) );
  nd02d0 U13380 ( .A1(n2678), .A2(n2677), .ZN(N8096) );
  aoi21d1 U13381 ( .B1(n1100), .B2(n1049), .A(n1139), .ZN(n2680) );
  nr04d0 U13382 ( .A1(n1341), .A2(n1308), .A3(n1255), .A4(n1206), .ZN(n2679)
         );
  oaim311d1 U13383 ( .C1(n977), .C2(n1110), .C3(n1014), .A(n2680), .B(n2679), 
        .ZN(N8085) );
  nr02d0 U13384 ( .A1(n1207), .A2(n1159), .ZN(n2683) );
  oai21d1 U13385 ( .B1(n1014), .B2(n1057), .A(n1103), .ZN(n2682) );
  nr03d0 U13386 ( .A1(n1251), .A2(n1346), .A3(n1300), .ZN(n2681) );
  nd03d0 U13387 ( .A1(n2683), .A2(n2682), .A3(n2681), .ZN(N8074) );
  nr02d0 U13388 ( .A1(n1026), .A2(n978), .ZN(n2686) );
  aoi21d1 U13389 ( .B1(n1101), .B2(n1049), .A(n1149), .ZN(n2685) );
  nr04d0 U13390 ( .A1(n1340), .A2(n1308), .A3(n1255), .A4(n1206), .ZN(n2684)
         );
  oai211d1 U13391 ( .C1(n2686), .C2(n1128), .A(n2685), .B(n2684), .ZN(N8064)
         );
  nr03d0 U13392 ( .A1(n1118), .A2(n1206), .A3(n1163), .ZN(n2688) );
  nr03d0 U13393 ( .A1(n1250), .A2(n1346), .A3(n1303), .ZN(n2687) );
  nd02d0 U13394 ( .A1(n2688), .A2(n2687), .ZN(N8054) );
  aoi311d1 U13395 ( .C1(n1001), .C2(n963), .C3(n1043), .A(n1137), .B(
        num_images[3]), .ZN(n2690) );
  nr04d0 U13396 ( .A1(n1340), .A2(n1308), .A3(n1229), .A4(n1206), .ZN(n2689)
         );
  nd02d0 U13397 ( .A1(n2690), .A2(n2689), .ZN(N8044) );
  aoi211d1 U13398 ( .C1(n1062), .C2(n1008), .A(n1145), .B(n1105), .ZN(n2692)
         );
  nr04d0 U13399 ( .A1(n1340), .A2(n1308), .A3(n1231), .A4(n1205), .ZN(n2691)
         );
  nd02d0 U13400 ( .A1(n2692), .A2(n2691), .ZN(N8034) );
  nr02d0 U13401 ( .A1(n1162), .A2(n1107), .ZN(n2695) );
  oai21d1 U13402 ( .B1(n1014), .B2(n968), .A(n1061), .ZN(n2694) );
  nr04d0 U13403 ( .A1(n1341), .A2(n1309), .A3(n1255), .A4(n1206), .ZN(n2693)
         );
  nd03d0 U13404 ( .A1(n2695), .A2(n2694), .A3(n2693), .ZN(N8025) );
  nr03d0 U13405 ( .A1(n1070), .A2(n1143), .A3(n1116), .ZN(n2697) );
  nr04d0 U13406 ( .A1(n1340), .A2(n1308), .A3(num_images[6]), .A4(n1206), .ZN(
        n2696) );
  nd02d0 U13407 ( .A1(n2697), .A2(n2696), .ZN(N8016) );
  aoi21d1 U13408 ( .B1(n1012), .B2(n964), .A(n1063), .ZN(n2700) );
  nr02d0 U13409 ( .A1(n1162), .A2(n1118), .ZN(n2699) );
  nr04d0 U13410 ( .A1(n1341), .A2(n1308), .A3(n1236), .A4(n1205), .ZN(n2698)
         );
  nd03d0 U13411 ( .A1(n2700), .A2(n2699), .A3(n2698), .ZN(N8008) );
  nr04d0 U13412 ( .A1(n1158), .A2(n1118), .A3(n1041), .A4(n1023), .ZN(n2702)
         );
  nr04d0 U13413 ( .A1(n1340), .A2(n1309), .A3(n1235), .A4(n1206), .ZN(n2701)
         );
  nd02d0 U13414 ( .A1(n2702), .A2(n2701), .ZN(N8001) );
  nr02d0 U13415 ( .A1(n1202), .A2(n1160), .ZN(n2705) );
  nr03d0 U13416 ( .A1(n1251), .A2(n1345), .A3(n1270), .ZN(n2704) );
  nr04d0 U13417 ( .A1(n1117), .A2(n1070), .A3(n1026), .A4(n979), .ZN(n2703) );
  nd03d0 U13418 ( .A1(n2705), .A2(n2704), .A3(n2703), .ZN(N7997) );
  or02d0 U13419 ( .A1(n506), .A2(n1219), .Z(n2714) );
  an02d0 U13420 ( .A1(n1114), .A2(n956), .Z(n2707) );
  nr03d0 U13421 ( .A1(n2707), .A2(n1071), .A3(n501), .ZN(n2706) );
  aoim21d1 U13422 ( .B1(n1092), .B2(n956), .A(n2706), .ZN(n2709) );
  aon211d1 U13423 ( .C1(n1047), .C2(n501), .B(n2707), .A(n2709), .ZN(n2708) );
  oai211d1 U13424 ( .C1(n504), .C2(n1133), .A(n2714), .B(n2708), .ZN(n2719) );
  aoim22d1 U13425 ( .A1(n961), .A2(n512), .B1(n1035), .B2(n500), .Z(n2710) );
  aoi211d1 U13426 ( .C1(n500), .C2(n1034), .A(n2721), .B(n2710), .ZN(n2718) );
  nd02d0 U13427 ( .A1(n1309), .A2(n418), .ZN(n2711) );
  oai21d1 U13428 ( .B1(N3180), .B2(n1267), .A(n2711), .ZN(n2717) );
  nd03d0 U13429 ( .A1(n2711), .A2(n1258), .A3(N3180), .ZN(n2712) );
  oai21d1 U13430 ( .B1(n1279), .B2(n418), .A(n2712), .ZN(n2713) );
  aoi321d1 U13431 ( .C1(n504), .C2(n1173), .C3(n2714), .B1(n1218), .B2(n506), 
        .A(n2713), .ZN(n2715) );
  aor21d1 U13432 ( .B1(n2717), .B2(n2722), .A(n2715), .Z(n2716) );
  oai321d1 U13433 ( .C1(n2719), .C2(n2718), .C3(n2717), .B1(n1343), .B2(n419), 
        .A(n2716), .ZN(n2720) );
  oaim21d1 U13434 ( .B1(n419), .B2(n1331), .A(n2720), .ZN(N4760) );
  or02d0 U13435 ( .A1(\lt_82/A[5] ), .A2(n1218), .Z(n2731) );
  an02d0 U13436 ( .A1(n1114), .A2(n2739), .Z(n2724) );
  nr03d0 U13437 ( .A1(n2724), .A2(n1071), .A3(n2784), .ZN(n2723) );
  aoim21d1 U13438 ( .B1(n1092), .B2(n2739), .A(n2723), .ZN(n2726) );
  aon211d1 U13439 ( .C1(n1047), .C2(n2784), .B(n2724), .A(n2726), .ZN(n2725)
         );
  oai211d1 U13440 ( .C1(\lt_82/A[4] ), .C2(n1164), .A(n2731), .B(n2725), .ZN(
        n2736) );
  aoim22d1 U13441 ( .A1(n961), .A2(n2741), .B1(n1035), .B2(count_image[1]), 
        .Z(n2727) );
  aoi211d1 U13442 ( .C1(count_image[1]), .C2(n1035), .A(n2740), .B(n2727), 
        .ZN(n2735) );
  nd02d0 U13443 ( .A1(n1309), .A2(n2742), .ZN(n2728) );
  oai21d1 U13444 ( .B1(count_image[6]), .B2(n1268), .A(n2728), .ZN(n2734) );
  nd03d0 U13445 ( .A1(n2728), .A2(n1269), .A3(count_image[6]), .ZN(n2729) );
  oai21d1 U13446 ( .B1(n1279), .B2(n2742), .A(n2729), .ZN(n2730) );
  aoi321d1 U13447 ( .C1(\lt_82/A[4] ), .C2(n1174), .C3(n2731), .B1(n1220), 
        .B2(\lt_82/A[5] ), .A(n2730), .ZN(n2732) );
  aor21d1 U13448 ( .B1(n2734), .B2(n2743), .A(n2732), .Z(n2733) );
  oai321d1 U13449 ( .C1(n2736), .C2(n2735), .C3(n2734), .B1(n1330), .B2(n2738), 
        .A(n2733), .ZN(n2737) );
  oaim21d1 U13450 ( .B1(n2738), .B2(n1331), .A(n2737), .ZN(N3187) );
  an02d1 U13451 ( .A1(N29403), .A2(N29404), .Z(n7615) );
  an02d1 U13452 ( .A1(N29399), .A2(N29400), .Z(n7621) );
  aoi22d1 U13454 ( .A1(reorder_A2[1]), .A2(n3594), .B1(N3877), .B2(n954), .ZN(
        n3591) );
  aoi22d1 U13455 ( .A1(reorder_A2[2]), .A2(n3594), .B1(N3878), .B2(n954), .ZN(
        n3595) );
  aoi22d1 U13456 ( .A1(reorder_A1[1]), .A2(n3623), .B1(N3877), .B2(n954), .ZN(
        n3624) );
  aoi22d1 U13457 ( .A1(reorder_A1[2]), .A2(n3623), .B1(N3878), .B2(n953), .ZN(
        n3626) );
  xr02d1 U13458 ( .A1(N29405), .A2(n7615), .Z(N4724) );
  xr02d1 U13459 ( .A1(N29404), .A2(N29403), .Z(N4723) );
  xr02d1 U13460 ( .A1(N29401), .A2(n7621), .Z(N3915) );
  xr02d1 U13461 ( .A1(N29400), .A2(N29399), .Z(N3914) );
endmodule


module controller_DW01_inc_0_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  ah01d1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ah01d1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ah01d1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ah01d1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ah01d1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ah01d1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ah01d1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  inv0d0 U1 ( .I(A[0]), .ZN(SUM[0]) );
  xr02d1 U2 ( .A1(carry[8]), .A2(A[8]), .Z(SUM[8]) );
endmodule


module controller ( clk, reset, start, image_buffer_valid, num_images, 
        finish_reordering, hash_calc_done, buffer_A1, buffer_I1, buffer_WEB1, 
        hash_A1, hash_A2, hash_I1, hash_WEB1, hash_WEB2, reorder_A1, 
        reorder_A2, reorder_WEB1, reorder_WEB2, controller_A1, controller_A2, 
        controller_I1, controller_I2, controller_WEB1, controller_WEB2, 
        controller_OEB1, controller_OEB2, controller_CSB1, controller_CSB2, 
        hash_start, reorder_start );
  input [8:0] num_images;
  input [11:0] buffer_A1;
  input [31:0] buffer_I1;
  input [11:0] hash_A1;
  input [11:0] hash_A2;
  input [31:0] hash_I1;
  input [11:0] reorder_A1;
  input [11:0] reorder_A2;
  output [11:0] controller_A1;
  output [11:0] controller_A2;
  output [31:0] controller_I1;
  output [31:0] controller_I2;
  input clk, reset, start, image_buffer_valid, finish_reordering,
         hash_calc_done, buffer_WEB1, hash_WEB1, hash_WEB2, reorder_WEB1,
         reorder_WEB2;
  output controller_WEB1, controller_WEB2, controller_OEB1, controller_OEB2,
         controller_CSB1, controller_CSB2, hash_start, reorder_start;
  wire   N23, N24, N25, N26, N27, N28, N29, N30, N31, N34, N38, N39, N40, N41,
         N42, N43, N44, N45, N46, N61, N62, N63, N64, N65, N66, N67, N68, N69,
         N70, N71, N72, n17, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n18, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73;
  wire   [1:0] current_state;
  wire   [8:0] current_image;
  wire   [1:0] next_state;
  wire   [8:0] next_image;
  assign controller_CSB2 = 1'b0;
  assign controller_CSB1 = 1'b0;
  assign controller_OEB2 = 1'b0;
  assign controller_OEB1 = 1'b0;
  assign controller_I2[0] = 1'b0;
  assign controller_I2[1] = 1'b0;
  assign controller_I2[2] = 1'b0;
  assign controller_I2[3] = 1'b0;
  assign controller_I2[4] = 1'b0;
  assign controller_I2[5] = 1'b0;
  assign controller_I2[6] = 1'b0;
  assign controller_I2[7] = 1'b0;
  assign controller_I2[8] = 1'b0;
  assign controller_I2[9] = 1'b0;
  assign controller_I2[10] = 1'b0;
  assign controller_I2[11] = 1'b0;
  assign controller_I2[12] = 1'b0;
  assign controller_I2[13] = 1'b0;
  assign controller_I2[14] = 1'b0;
  assign controller_I2[15] = 1'b0;
  assign controller_I2[16] = 1'b0;
  assign controller_I2[17] = 1'b0;
  assign controller_I2[18] = 1'b0;
  assign controller_I2[19] = 1'b0;
  assign controller_I2[20] = 1'b0;
  assign controller_I2[21] = 1'b0;
  assign controller_I2[22] = 1'b0;
  assign controller_I2[23] = 1'b0;
  assign controller_I2[24] = 1'b0;
  assign controller_I2[25] = 1'b0;
  assign controller_I2[26] = 1'b0;
  assign controller_I2[27] = 1'b0;
  assign controller_I2[28] = 1'b0;
  assign controller_I2[29] = 1'b0;
  assign controller_I2[30] = 1'b0;
  assign controller_I2[31] = 1'b0;

  lanhq1 \next_image_reg[0]  ( .E(N61), .D(N62), .Q(next_image[0]) );
  lanhq1 \next_image_reg[8]  ( .E(N61), .D(N70), .Q(next_image[8]) );
  lanhq1 \next_state_reg[0]  ( .E(N61), .D(N71), .Q(next_state[0]) );
  lanhq1 \next_state_reg[1]  ( .E(N61), .D(N72), .Q(next_state[1]) );
  lanhq1 \next_image_reg[7]  ( .E(N61), .D(N69), .Q(next_image[7]) );
  lanhq1 \next_image_reg[6]  ( .E(N61), .D(N68), .Q(next_image[6]) );
  lanhq1 \next_image_reg[5]  ( .E(N61), .D(N67), .Q(next_image[5]) );
  lanhq1 \next_image_reg[4]  ( .E(N61), .D(N66), .Q(next_image[4]) );
  lanhq1 \next_image_reg[3]  ( .E(N61), .D(N65), .Q(next_image[3]) );
  lanhq1 \next_image_reg[2]  ( .E(N61), .D(N64), .Q(next_image[2]) );
  lanhq1 \next_image_reg[1]  ( .E(N61), .D(N63), .Q(next_image[1]) );
  nd04d1 U13 ( .A1(n28), .A2(n24), .A3(n19), .A4(n71), .ZN(N61) );
  aoi22d1 U26 ( .A1(reorder_WEB2), .A2(n70), .B1(hash_WEB2), .B2(hash_start), 
        .ZN(n17) );
  aor222d1 U27 ( .A1(hash_WEB1), .A2(n14), .B1(reorder_WEB1), .B2(n70), .C1(
        buffer_WEB1), .C2(n6), .Z(controller_WEB1) );
  aor22d1 U28 ( .A1(buffer_I1[9]), .A2(n6), .B1(hash_I1[9]), .B2(n3), .Z(
        controller_I1[9]) );
  aor22d1 U29 ( .A1(buffer_I1[8]), .A2(n6), .B1(hash_I1[8]), .B2(n4), .Z(
        controller_I1[8]) );
  aor22d1 U30 ( .A1(buffer_I1[7]), .A2(n6), .B1(hash_I1[7]), .B2(n4), .Z(
        controller_I1[7]) );
  aor22d1 U31 ( .A1(buffer_I1[6]), .A2(n6), .B1(hash_I1[6]), .B2(n3), .Z(
        controller_I1[6]) );
  aor22d1 U32 ( .A1(buffer_I1[5]), .A2(n7), .B1(hash_I1[5]), .B2(n4), .Z(
        controller_I1[5]) );
  aor22d1 U33 ( .A1(buffer_I1[4]), .A2(n7), .B1(hash_I1[4]), .B2(n3), .Z(
        controller_I1[4]) );
  aor22d1 U34 ( .A1(buffer_I1[3]), .A2(n7), .B1(hash_I1[3]), .B2(n4), .Z(
        controller_I1[3]) );
  aor22d1 U35 ( .A1(buffer_I1[31]), .A2(n7), .B1(hash_I1[31]), .B2(n3), .Z(
        controller_I1[31]) );
  aor22d1 U36 ( .A1(buffer_I1[30]), .A2(n7), .B1(hash_I1[30]), .B2(n4), .Z(
        controller_I1[30]) );
  aor22d1 U37 ( .A1(buffer_I1[2]), .A2(n8), .B1(hash_I1[2]), .B2(n3), .Z(
        controller_I1[2]) );
  aor22d1 U38 ( .A1(buffer_I1[29]), .A2(n7), .B1(hash_I1[29]), .B2(n4), .Z(
        controller_I1[29]) );
  aor22d1 U39 ( .A1(buffer_I1[28]), .A2(n7), .B1(hash_I1[28]), .B2(n3), .Z(
        controller_I1[28]) );
  aor22d1 U40 ( .A1(buffer_I1[27]), .A2(n7), .B1(hash_I1[27]), .B2(n4), .Z(
        controller_I1[27]) );
  aor22d1 U41 ( .A1(buffer_I1[26]), .A2(n7), .B1(hash_I1[26]), .B2(n3), .Z(
        controller_I1[26]) );
  aor22d1 U42 ( .A1(buffer_I1[25]), .A2(n7), .B1(hash_I1[25]), .B2(n3), .Z(
        controller_I1[25]) );
  aor22d1 U43 ( .A1(buffer_I1[24]), .A2(n8), .B1(hash_I1[24]), .B2(n3), .Z(
        controller_I1[24]) );
  aor22d1 U44 ( .A1(buffer_I1[23]), .A2(n8), .B1(hash_I1[23]), .B2(n4), .Z(
        controller_I1[23]) );
  aor22d1 U45 ( .A1(buffer_I1[22]), .A2(n8), .B1(hash_I1[22]), .B2(n3), .Z(
        controller_I1[22]) );
  aor22d1 U46 ( .A1(buffer_I1[21]), .A2(n8), .B1(hash_I1[21]), .B2(n4), .Z(
        controller_I1[21]) );
  aor22d1 U47 ( .A1(buffer_I1[20]), .A2(n8), .B1(hash_I1[20]), .B2(n3), .Z(
        controller_I1[20]) );
  aor22d1 U48 ( .A1(buffer_I1[1]), .A2(n8), .B1(hash_I1[1]), .B2(n4), .Z(
        controller_I1[1]) );
  aor22d1 U49 ( .A1(buffer_I1[19]), .A2(n8), .B1(hash_I1[19]), .B2(n3), .Z(
        controller_I1[19]) );
  aor22d1 U50 ( .A1(buffer_I1[18]), .A2(n8), .B1(hash_I1[18]), .B2(n4), .Z(
        controller_I1[18]) );
  aor22d1 U51 ( .A1(buffer_I1[17]), .A2(n8), .B1(hash_I1[17]), .B2(n3), .Z(
        controller_I1[17]) );
  aor22d1 U52 ( .A1(buffer_I1[16]), .A2(n9), .B1(hash_I1[16]), .B2(n4), .Z(
        controller_I1[16]) );
  aor22d1 U53 ( .A1(buffer_I1[15]), .A2(n9), .B1(hash_I1[15]), .B2(n3), .Z(
        controller_I1[15]) );
  aor22d1 U54 ( .A1(buffer_I1[14]), .A2(n9), .B1(hash_I1[14]), .B2(n4), .Z(
        controller_I1[14]) );
  aor22d1 U55 ( .A1(buffer_I1[13]), .A2(n9), .B1(hash_I1[13]), .B2(hash_start), 
        .Z(controller_I1[13]) );
  aor22d1 U56 ( .A1(buffer_I1[12]), .A2(n9), .B1(hash_I1[12]), .B2(n14), .Z(
        controller_I1[12]) );
  aor22d1 U57 ( .A1(buffer_I1[11]), .A2(n9), .B1(hash_I1[11]), .B2(n3), .Z(
        controller_I1[11]) );
  aor22d1 U58 ( .A1(buffer_I1[10]), .A2(n9), .B1(hash_I1[10]), .B2(n4), .Z(
        controller_I1[10]) );
  aor22d1 U59 ( .A1(buffer_I1[0]), .A2(n6), .B1(hash_I1[0]), .B2(n14), .Z(
        controller_I1[0]) );
  aor22d1 U60 ( .A1(hash_A2[9]), .A2(n14), .B1(reorder_A2[9]), .B2(n13), .Z(
        controller_A2[9]) );
  aor22d1 U61 ( .A1(hash_A2[8]), .A2(n14), .B1(reorder_A2[8]), .B2(n13), .Z(
        controller_A2[8]) );
  aor22d1 U62 ( .A1(hash_A2[7]), .A2(n14), .B1(reorder_A2[7]), .B2(n13), .Z(
        controller_A2[7]) );
  aor22d1 U63 ( .A1(hash_A2[6]), .A2(n14), .B1(reorder_A2[6]), .B2(n70), .Z(
        controller_A2[6]) );
  aor22d1 U64 ( .A1(hash_A2[5]), .A2(n14), .B1(reorder_A2[5]), .B2(n13), .Z(
        controller_A2[5]) );
  aor22d1 U65 ( .A1(hash_A2[4]), .A2(n14), .B1(reorder_A2[4]), .B2(n13), .Z(
        controller_A2[4]) );
  aor22d1 U66 ( .A1(hash_A2[3]), .A2(n14), .B1(reorder_A2[3]), .B2(n13), .Z(
        controller_A2[3]) );
  aor22d1 U67 ( .A1(hash_A2[2]), .A2(n14), .B1(reorder_A2[2]), .B2(n13), .Z(
        controller_A2[2]) );
  aor22d1 U68 ( .A1(hash_A2[1]), .A2(n14), .B1(reorder_A2[1]), .B2(n70), .Z(
        controller_A2[1]) );
  aor22d1 U69 ( .A1(hash_A2[11]), .A2(n14), .B1(reorder_A2[11]), .B2(n70), .Z(
        controller_A2[11]) );
  aor22d1 U70 ( .A1(hash_A2[10]), .A2(n14), .B1(reorder_A2[10]), .B2(n70), .Z(
        controller_A2[10]) );
  aor22d1 U71 ( .A1(hash_A2[0]), .A2(n14), .B1(reorder_A2[0]), .B2(n70), .Z(
        controller_A2[0]) );
  aor222d1 U72 ( .A1(hash_A1[9]), .A2(n4), .B1(reorder_A1[9]), .B2(n13), .C1(
        buffer_A1[9]), .C2(n6), .Z(controller_A1[9]) );
  aor222d1 U73 ( .A1(hash_A1[8]), .A2(n3), .B1(reorder_A1[8]), .B2(
        reorder_start), .C1(buffer_A1[8]), .C2(n6), .Z(controller_A1[8]) );
  aor222d1 U74 ( .A1(hash_A1[7]), .A2(n3), .B1(reorder_A1[7]), .B2(
        reorder_start), .C1(buffer_A1[7]), .C2(n6), .Z(controller_A1[7]) );
  aor222d1 U75 ( .A1(hash_A1[6]), .A2(n4), .B1(reorder_A1[6]), .B2(
        reorder_start), .C1(buffer_A1[6]), .C2(n5), .Z(controller_A1[6]) );
  aor222d1 U76 ( .A1(hash_A1[5]), .A2(n3), .B1(reorder_A1[5]), .B2(
        reorder_start), .C1(buffer_A1[5]), .C2(n5), .Z(controller_A1[5]) );
  aor222d1 U77 ( .A1(hash_A1[4]), .A2(n3), .B1(reorder_A1[4]), .B2(
        reorder_start), .C1(buffer_A1[4]), .C2(n5), .Z(controller_A1[4]) );
  aor222d1 U78 ( .A1(hash_A1[3]), .A2(n4), .B1(reorder_A1[3]), .B2(
        reorder_start), .C1(buffer_A1[3]), .C2(n5), .Z(controller_A1[3]) );
  aor222d1 U79 ( .A1(hash_A1[2]), .A2(n4), .B1(reorder_A1[2]), .B2(
        reorder_start), .C1(buffer_A1[2]), .C2(n5), .Z(controller_A1[2]) );
  aor222d1 U80 ( .A1(hash_A1[1]), .A2(n3), .B1(reorder_A1[1]), .B2(n70), .C1(
        buffer_A1[1]), .C2(n5), .Z(controller_A1[1]) );
  aor222d1 U81 ( .A1(hash_A1[11]), .A2(n4), .B1(reorder_A1[11]), .B2(n70), 
        .C1(buffer_A1[11]), .C2(n5), .Z(controller_A1[11]) );
  aor222d1 U82 ( .A1(hash_A1[10]), .A2(n3), .B1(reorder_A1[10]), .B2(n13), 
        .C1(buffer_A1[10]), .C2(n5), .Z(controller_A1[10]) );
  aor222d1 U83 ( .A1(hash_A1[0]), .A2(n4), .B1(reorder_A1[0]), .B2(n70), .C1(
        buffer_A1[0]), .C2(n5), .Z(controller_A1[0]) );
  oai211d1 U84 ( .C1(n67), .C2(n69), .A(n20), .B(n21), .ZN(N71) );
  aoi22d1 U85 ( .A1(n22), .A2(N34), .B1(start), .B2(n23), .ZN(n21) );
  oai22d1 U86 ( .A1(finish_reordering), .A2(n19), .B1(n26), .B2(n24), .ZN(n25)
         );
  aor22d1 U87 ( .A1(current_image[8]), .A2(n27), .B1(N46), .B2(n66), .Z(N70)
         );
  aor22d1 U88 ( .A1(current_image[7]), .A2(n27), .B1(N45), .B2(n66), .Z(N69)
         );
  aor22d1 U89 ( .A1(current_image[6]), .A2(n27), .B1(N44), .B2(n66), .Z(N68)
         );
  aor22d1 U90 ( .A1(current_image[5]), .A2(n27), .B1(N43), .B2(n66), .Z(N67)
         );
  aor22d1 U91 ( .A1(current_image[4]), .A2(n27), .B1(N42), .B2(n66), .Z(N66)
         );
  aor22d1 U92 ( .A1(current_image[3]), .A2(n27), .B1(N41), .B2(n66), .Z(N65)
         );
  aor22d1 U93 ( .A1(current_image[2]), .A2(n27), .B1(N40), .B2(n66), .Z(N64)
         );
  aor22d1 U94 ( .A1(current_image[1]), .A2(n27), .B1(N39), .B2(n66), .Z(N63)
         );
  aor22d1 U95 ( .A1(current_image[0]), .A2(n27), .B1(N38), .B2(n66), .Z(N62)
         );
  controller_DW01_inc_0_DW01_inc_1 add_104 ( .A(current_image), .SUM({N46, N45, 
        N44, N43, N42, N41, N40, N39, N38}) );
  dfcrq1 \current_image_reg[8]  ( .D(next_image[8]), .CP(clk), .CDN(n73), .Q(
        current_image[8]) );
  dfcrq1 \current_image_reg[7]  ( .D(next_image[7]), .CP(clk), .CDN(n73), .Q(
        current_image[7]) );
  dfcrq1 \current_image_reg[6]  ( .D(next_image[6]), .CP(clk), .CDN(n73), .Q(
        current_image[6]) );
  dfcrq1 \current_image_reg[3]  ( .D(next_image[3]), .CP(clk), .CDN(n73), .Q(
        current_image[3]) );
  dfcrq1 \current_image_reg[2]  ( .D(next_image[2]), .CP(clk), .CDN(n73), .Q(
        current_image[2]) );
  dfcrq1 \current_image_reg[4]  ( .D(next_image[4]), .CP(clk), .CDN(n73), .Q(
        current_image[4]) );
  dfcrq1 \current_image_reg[5]  ( .D(next_image[5]), .CP(clk), .CDN(n73), .Q(
        current_image[5]) );
  dfcrq1 \current_image_reg[1]  ( .D(next_image[1]), .CP(clk), .CDN(n73), .Q(
        current_image[1]) );
  dfcrq1 \current_image_reg[0]  ( .D(next_image[0]), .CP(clk), .CDN(n73), .Q(
        current_image[0]) );
  dfcrq1 \current_state_reg[1]  ( .D(next_state[1]), .CP(clk), .CDN(n73), .Q(
        current_state[1]) );
  dfcrq1 \current_state_reg[0]  ( .D(next_state[0]), .CP(clk), .CDN(n73), .Q(
        current_state[0]) );
  buffd1 U3 ( .I(n13), .Z(reorder_start) );
  inv0d1 U4 ( .I(n24), .ZN(n3) );
  inv0d1 U5 ( .I(n24), .ZN(n4) );
  inv0d0 U6 ( .I(n10), .ZN(n5) );
  buffd1 U7 ( .I(hash_start), .Z(n14) );
  inv0d0 U8 ( .I(n20), .ZN(n66) );
  buffd1 U9 ( .I(n2), .Z(n10) );
  inv0d0 U10 ( .I(n11), .ZN(n6) );
  buffd1 U11 ( .I(n2), .Z(n11) );
  inv0d0 U12 ( .I(n24), .ZN(hash_start) );
  inv0d0 U14 ( .I(n19), .ZN(n13) );
  inv0d0 U15 ( .I(n19), .ZN(n70) );
  inv0d0 U16 ( .I(n12), .ZN(n7) );
  inv0d0 U17 ( .I(n12), .ZN(n8) );
  buffd1 U18 ( .I(n2), .Z(n12) );
  inv0d0 U19 ( .I(n23), .ZN(n71) );
  inv0d0 U20 ( .I(n39), .ZN(n63) );
  nd04d1 U21 ( .A1(n26), .A2(n10), .A3(n19), .A4(n71), .ZN(n27) );
  nd02d1 U22 ( .A1(n26), .A2(n4), .ZN(n20) );
  inv0d0 U23 ( .I(n33), .ZN(n35) );
  nd02d1 U24 ( .A1(n67), .A2(n10), .ZN(N72) );
  inv0d0 U25 ( .I(n50), .ZN(n61) );
  inv0d0 U96 ( .I(n11), .ZN(n9) );
  inv0d0 U97 ( .I(n16), .ZN(n15) );
  or02d0 U98 ( .A1(n69), .A2(current_state[1]), .Z(n2) );
  inv0d0 U99 ( .I(current_state[0]), .ZN(n69) );
  nd03d1 U100 ( .A1(n10), .A2(n71), .A3(n17), .ZN(controller_WEB2) );
  nd02d1 U101 ( .A1(current_state[1]), .A2(n69), .ZN(n24) );
  nd02d1 U102 ( .A1(current_state[1]), .A2(current_state[0]), .ZN(n19) );
  nr02d1 U103 ( .A1(current_state[0]), .A2(current_state[1]), .ZN(n23) );
  nd02d1 U104 ( .A1(image_buffer_valid), .A2(n72), .ZN(n28) );
  inv0d1 U105 ( .I(reset), .ZN(n73) );
  an12d1 U106 ( .A2(hash_calc_done), .A1(n54), .Z(n26) );
  nr02d1 U107 ( .A1(n24), .A2(n72), .ZN(n22) );
  inv0d0 U108 ( .I(N23), .ZN(n55) );
  inv0d0 U109 ( .I(n34), .ZN(N30) );
  inv0d0 U110 ( .I(n25), .ZN(n67) );
  inv0d0 U111 ( .I(hash_calc_done), .ZN(n72) );
  inv0d0 U112 ( .I(N27), .ZN(n57) );
  inv0d0 U113 ( .I(current_image[8]), .ZN(n65) );
  inv0d0 U114 ( .I(N26), .ZN(n56) );
  inv0d0 U115 ( .I(current_image[1]), .ZN(n58) );
  inv0d0 U116 ( .I(current_image[2]), .ZN(n59) );
  inv0d0 U117 ( .I(current_image[6]), .ZN(n62) );
  inv0d0 U118 ( .I(current_image[3]), .ZN(n60) );
  inv0d0 U119 ( .I(current_image[7]), .ZN(n64) );
  inv0d0 U120 ( .I(num_images[0]), .ZN(n16) );
  nd12d0 U121 ( .A1(num_images[1]), .A2(n16), .ZN(n18) );
  oaim21d1 U122 ( .B1(n15), .B2(num_images[1]), .A(n18), .ZN(N23) );
  or02d0 U123 ( .A1(n18), .A2(num_images[2]), .Z(n29) );
  oaim21d1 U124 ( .B1(n18), .B2(num_images[2]), .A(n29), .ZN(N24) );
  or02d0 U125 ( .A1(n29), .A2(num_images[3]), .Z(n30) );
  oaim21d1 U126 ( .B1(n29), .B2(num_images[3]), .A(n30), .ZN(N25) );
  or02d0 U127 ( .A1(n30), .A2(num_images[4]), .Z(n31) );
  oaim21d1 U128 ( .B1(n30), .B2(num_images[4]), .A(n31), .ZN(N26) );
  or02d0 U129 ( .A1(n31), .A2(num_images[5]), .Z(n32) );
  oaim21d1 U130 ( .B1(n31), .B2(num_images[5]), .A(n32), .ZN(N27) );
  nr02d0 U131 ( .A1(n32), .A2(num_images[6]), .ZN(n33) );
  oaim21d1 U132 ( .B1(n32), .B2(num_images[6]), .A(n35), .ZN(N28) );
  xr02d1 U133 ( .A1(num_images[7]), .A2(n33), .Z(N29) );
  nr03d0 U134 ( .A1(num_images[7]), .A2(num_images[8]), .A3(n35), .ZN(N31) );
  oan211d1 U135 ( .C1(n35), .C2(num_images[7]), .B(num_images[8]), .A(N31), 
        .ZN(n34) );
  an02d0 U136 ( .A1(current_image[0]), .A2(n15), .Z(n36) );
  oai22d1 U137 ( .A1(current_image[1]), .A2(n36), .B1(n36), .B2(n55), .ZN(n38)
         );
  nr02d0 U138 ( .A1(n62), .A2(N28), .ZN(n39) );
  nr02d0 U139 ( .A1(n64), .A2(N29), .ZN(n46) );
  nr02d0 U140 ( .A1(n39), .A2(n46), .ZN(n37) );
  oai211d1 U141 ( .C1(N30), .C2(n65), .A(n38), .B(n37), .ZN(n53) );
  nr02d0 U142 ( .A1(n60), .A2(N25), .ZN(n49) );
  or02d0 U143 ( .A1(N24), .A2(n59), .Z(n48) );
  nd02d0 U144 ( .A1(current_image[5]), .A2(n57), .ZN(n50) );
  nr02d0 U145 ( .A1(n15), .A2(current_image[0]), .ZN(n41) );
  aon211d1 U146 ( .C1(n41), .C2(n58), .B(N23), .A(n48), .ZN(n40) );
  aoim21d1 U147 ( .B1(n58), .B2(n41), .A(n40), .ZN(n42) );
  aoi221d1 U148 ( .B1(N25), .B2(n60), .C1(N24), .C2(n59), .A(n42), .ZN(n43) );
  an02d0 U149 ( .A1(current_image[4]), .A2(n56), .Z(n51) );
  oai322d1 U150 ( .C1(n43), .C2(n49), .C3(n51), .A1(current_image[4]), .A2(n56), .B1(current_image[5]), .B2(n57), .ZN(n44) );
  aoi322d1 U151 ( .C1(n63), .C2(n50), .C3(n44), .A1(N29), .A2(n64), .B1(N28), 
        .B2(n62), .ZN(n45) );
  aoim211d1 U152 ( .C1(n65), .C2(N30), .A(n46), .B(n45), .ZN(n47) );
  aoi211d1 U153 ( .C1(N30), .C2(n65), .A(N31), .B(n47), .ZN(n54) );
  nd13d1 U154 ( .A1(n49), .A2(n48), .A3(n54), .ZN(n52) );
  nr04d0 U155 ( .A1(n53), .A2(n52), .A3(n51), .A4(n61), .ZN(N34) );
endmodule


module top_syn ( clk, reset, pixel_data, pixel_valid, start, num_images, 
        image_header, image_buffer_valid, hash_calc_done, finish_reordering, 
        temp_new_reference, new_reference_is_done, last_image, count_image );
  input [7:0] pixel_data;
  input [8:0] num_images;
  input [8:0] image_header;
  output [8:0] temp_new_reference;
  output [8:0] last_image;
  output [8:0] count_image;
  input clk, reset, pixel_valid, start;
  output image_buffer_valid, hash_calc_done, finish_reordering,
         new_reference_is_done;
  wire   hash_start, reorder_start, WEB1, WEB2, n1;
  wire   [15:0] sum;
  wire   [31:0] buffer_I1;
  wire   [11:0] buffer_A1;
  wire   [11:0] hash_A1;
  wire   [11:0] hash_A2;
  wire   [31:0] O2;
  wire   [31:0] hash_I1;
  wire   [11:0] reorder_A1;
  wire   [11:0] reorder_A2;
  wire   [31:0] O1;
  wire   [31:0] I1;
  wire   [31:0] I2;
  wire   [11:0] A1;
  wire   [11:0] A2;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26;

  dpram4096x32_CB RAM_U1 ( .A1(A1), .I1(I1), .O1(O1), .A2(A2), .I2({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .O2(O2), .CEB1(clk), .CEB2(clk), 
        .OEB1(1'b0), .CSB1(1'b0), .WEB1(WEB1), .OEB2(1'b0), .CSB2(1'b0), 
        .WEB2(WEB2) );
  image_buffer u_image_buffer ( .clk(clk), .reset(reset), .pixel_data(
        pixel_data), .pixel_valid(pixel_valid), .image_buffer_valid(
        image_buffer_valid), .sum(sum), .buffer_I1({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, buffer_I1[7:0]}), .buffer_A1(buffer_A1) );
  hash_calc u_hash_calc ( .clk(clk), .reset(reset), .image_header(image_header), .hash_start(hash_start), .sum(sum), .hash_calc_done(hash_calc_done), 
        .hash_O2(O2), .hash_I1(hash_I1), .hash_A1(hash_A1), .hash_A2({
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, hash_A2[8:0]}) );
  reordering u_reordering ( .clk(clk), .reset(reset), .num_images(num_images), 
        .reorder_start(n1), .temp_new_reference(temp_new_reference), 
        .new_reference_is_done(new_reference_is_done), .count_image(
        count_image), .last_image(last_image), .finish_reordering(
        finish_reordering), .reorder_O1(O1), .reorder_O2(O2), .reorder_A1(
        reorder_A1), .reorder_A2(reorder_A2) );
  controller u_controller ( .clk(clk), .reset(reset), .start(start), 
        .image_buffer_valid(image_buffer_valid), .num_images(num_images), 
        .finish_reordering(finish_reordering), .hash_calc_done(hash_calc_done), 
        .buffer_A1(buffer_A1), .buffer_I1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, buffer_I1[7:0]}), .buffer_WEB1(
        1'b0), .hash_A1(hash_A1), .hash_A2({1'b0, 1'b0, 1'b0, hash_A2[8:0]}), 
        .hash_I1(hash_I1), .hash_WEB1(1'b0), .hash_WEB2(1'b1), .reorder_A1(
        reorder_A1), .reorder_A2(reorder_A2), .reorder_WEB1(1'b1), 
        .reorder_WEB2(1'b1), .controller_A1(A1), .controller_A2(A2), 
        .controller_I1(I1), .controller_WEB1(WEB1), .controller_WEB2(WEB2), 
        .hash_start(hash_start), .reorder_start(reorder_start) );
  buffd1 U1 ( .I(reorder_start), .Z(n1) );
endmodule

module dpram4096x32_CB(A1, A2, CEB1, CEB2, WEB1, WEB2, OEB1, OEB2, CSB1, CSB2, I1, I2, O1, O2);
	input [11:0] A1;
	input CEB1,WEB1, OEB1, CSB1;
	input [31:0] I1;
	output [31:0] O1;
	input [11:0] A2;
	input CEB2,WEB2, OEB2, CSB2;
	input [31:0] I2;
	output [31:0] O2;
endmodule



